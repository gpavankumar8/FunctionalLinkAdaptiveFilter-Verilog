`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author: Pavan Kumar
// Create Date: 29-07-2024
// Module name: log_sin_cos_LUT_10QP.v
// The first and last entry after/before Inf in logsin and logcos has been set to -8 due to 4.12 limitations
//////////////////////////////////////////////////////////////////////////////////

module log_sin_cos_LUT_10QP
(
    input      [ 9:0] x_in1, x_in2, x_in3,
    output reg [15:0] logsin1, logsin2, logsin3, logcos1, logcos2, logcos3
);

    wire [15:0] mux_in_cos0, mux_in_sin0, mux_in_cos1, mux_in_sin1, mux_in_cos2, mux_in_sin2, mux_in_cos3, mux_in_sin3, mux_in_cos4, mux_in_sin4, mux_in_cos5, mux_in_sin5, mux_in_cos6, mux_in_sin6, mux_in_cos7, mux_in_sin7, mux_in_cos8, mux_in_sin8, mux_in_cos9, mux_in_sin9, mux_in_cos10, mux_in_sin10, mux_in_cos11, mux_in_sin11, mux_in_cos12, mux_in_sin12, mux_in_cos13, mux_in_sin13, mux_in_cos14, mux_in_sin14, mux_in_cos15, mux_in_sin15, mux_in_cos16, mux_in_sin16, mux_in_cos17, mux_in_sin17, mux_in_cos18, mux_in_sin18, mux_in_cos19, mux_in_sin19, mux_in_cos20, mux_in_sin20, mux_in_cos21, mux_in_sin21, mux_in_cos22, mux_in_sin22, mux_in_cos23, mux_in_sin23, mux_in_cos24, mux_in_sin24, mux_in_cos25, mux_in_sin25, mux_in_cos26, mux_in_sin26, mux_in_cos27, mux_in_sin27, mux_in_cos28, mux_in_sin28, mux_in_cos29, mux_in_sin29, mux_in_cos30, mux_in_sin30, mux_in_cos31, mux_in_sin31, mux_in_cos32, mux_in_sin32, mux_in_cos33, mux_in_sin33, mux_in_cos34, mux_in_sin34, mux_in_cos35, mux_in_sin35, mux_in_cos36, mux_in_sin36, mux_in_cos37, mux_in_sin37, mux_in_cos38, mux_in_sin38, mux_in_cos39, mux_in_sin39, mux_in_cos40, mux_in_sin40, mux_in_cos41, mux_in_sin41, mux_in_cos42, mux_in_sin42, mux_in_cos43, mux_in_sin43, mux_in_cos44, mux_in_sin44, mux_in_cos45, mux_in_sin45, mux_in_cos46, mux_in_sin46, mux_in_cos47, mux_in_sin47, mux_in_cos48, mux_in_sin48, mux_in_cos49, mux_in_sin49, mux_in_cos50, mux_in_sin50, mux_in_cos51, mux_in_sin51, mux_in_cos52, mux_in_sin52, mux_in_cos53, mux_in_sin53, mux_in_cos54, mux_in_sin54, mux_in_cos55, mux_in_sin55, mux_in_cos56, mux_in_sin56, mux_in_cos57, mux_in_sin57, mux_in_cos58, mux_in_sin58, mux_in_cos59, mux_in_sin59, mux_in_cos60, mux_in_sin60, mux_in_cos61, mux_in_sin61, mux_in_cos62, mux_in_sin62, mux_in_cos63, mux_in_sin63, mux_in_cos64, mux_in_sin64, mux_in_cos65, mux_in_sin65, mux_in_cos66, mux_in_sin66, mux_in_cos67, mux_in_sin67, mux_in_cos68, mux_in_sin68, mux_in_cos69, mux_in_sin69, mux_in_cos70, mux_in_sin70, mux_in_cos71, mux_in_sin71, mux_in_cos72, mux_in_sin72, mux_in_cos73, mux_in_sin73, mux_in_cos74, mux_in_sin74, mux_in_cos75, mux_in_sin75, mux_in_cos76, mux_in_sin76, mux_in_cos77, mux_in_sin77, mux_in_cos78, mux_in_sin78, mux_in_cos79, mux_in_sin79, mux_in_cos80, mux_in_sin80, mux_in_cos81, mux_in_sin81, mux_in_cos82, mux_in_sin82, mux_in_cos83, mux_in_sin83, mux_in_cos84, mux_in_sin84, mux_in_cos85, mux_in_sin85, mux_in_cos86, mux_in_sin86, mux_in_cos87, mux_in_sin87, mux_in_cos88, mux_in_sin88, mux_in_cos89, mux_in_sin89, mux_in_cos90, mux_in_sin90, mux_in_cos91, mux_in_sin91, mux_in_cos92, mux_in_sin92, mux_in_cos93, mux_in_sin93, mux_in_cos94, mux_in_sin94, mux_in_cos95, mux_in_sin95, mux_in_cos96, mux_in_sin96, mux_in_cos97, mux_in_sin97, mux_in_cos98, mux_in_sin98, mux_in_cos99, mux_in_sin99, mux_in_cos100, mux_in_sin100, mux_in_cos101, mux_in_sin101, mux_in_cos102, mux_in_sin102, mux_in_cos103, mux_in_sin103, mux_in_cos104, mux_in_sin104, mux_in_cos105, mux_in_sin105, mux_in_cos106, mux_in_sin106, mux_in_cos107, mux_in_sin107, mux_in_cos108, mux_in_sin108, mux_in_cos109, mux_in_sin109, mux_in_cos110, mux_in_sin110, mux_in_cos111, mux_in_sin111, mux_in_cos112, mux_in_sin112, mux_in_cos113, mux_in_sin113, mux_in_cos114, mux_in_sin114, mux_in_cos115, mux_in_sin115, mux_in_cos116, mux_in_sin116, mux_in_cos117, mux_in_sin117, mux_in_cos118, mux_in_sin118, mux_in_cos119, mux_in_sin119, mux_in_cos120, mux_in_sin120, mux_in_cos121, mux_in_sin121, mux_in_cos122, mux_in_sin122, mux_in_cos123, mux_in_sin123, mux_in_cos124, mux_in_sin124, mux_in_cos125, mux_in_sin125, mux_in_cos126, mux_in_sin126, mux_in_cos127, mux_in_sin127, mux_in_cos128, mux_in_sin128, mux_in_cos129, mux_in_sin129, mux_in_cos130, mux_in_sin130, mux_in_cos131, mux_in_sin131, mux_in_cos132, mux_in_sin132, mux_in_cos133, mux_in_sin133, mux_in_cos134, mux_in_sin134, mux_in_cos135, mux_in_sin135, mux_in_cos136, mux_in_sin136, mux_in_cos137, mux_in_sin137, mux_in_cos138, mux_in_sin138, mux_in_cos139, mux_in_sin139, mux_in_cos140, mux_in_sin140, mux_in_cos141, mux_in_sin141, mux_in_cos142, mux_in_sin142, mux_in_cos143, mux_in_sin143, mux_in_cos144, mux_in_sin144, mux_in_cos145, mux_in_sin145, mux_in_cos146, mux_in_sin146, mux_in_cos147, mux_in_sin147, mux_in_cos148, mux_in_sin148, mux_in_cos149, mux_in_sin149, mux_in_cos150, mux_in_sin150, mux_in_cos151, mux_in_sin151, mux_in_cos152, mux_in_sin152, mux_in_cos153, mux_in_sin153, mux_in_cos154, mux_in_sin154, mux_in_cos155, mux_in_sin155, mux_in_cos156, mux_in_sin156, mux_in_cos157, mux_in_sin157, mux_in_cos158, mux_in_sin158, mux_in_cos159, mux_in_sin159, mux_in_cos160, mux_in_sin160, mux_in_cos161, mux_in_sin161, mux_in_cos162, mux_in_sin162, mux_in_cos163, mux_in_sin163, mux_in_cos164, mux_in_sin164, mux_in_cos165, mux_in_sin165, mux_in_cos166, mux_in_sin166, mux_in_cos167, mux_in_sin167, mux_in_cos168, mux_in_sin168, mux_in_cos169, mux_in_sin169, mux_in_cos170, mux_in_sin170, mux_in_cos171, mux_in_sin171, mux_in_cos172, mux_in_sin172, mux_in_cos173, mux_in_sin173, mux_in_cos174, mux_in_sin174, mux_in_cos175, mux_in_sin175, mux_in_cos176, mux_in_sin176, mux_in_cos177, mux_in_sin177, mux_in_cos178, mux_in_sin178, mux_in_cos179, mux_in_sin179, mux_in_cos180, mux_in_sin180, mux_in_cos181, mux_in_sin181, mux_in_cos182, mux_in_sin182, mux_in_cos183, mux_in_sin183, mux_in_cos184, mux_in_sin184, mux_in_cos185, mux_in_sin185, mux_in_cos186, mux_in_sin186, mux_in_cos187, mux_in_sin187, mux_in_cos188, mux_in_sin188, mux_in_cos189, mux_in_sin189, mux_in_cos190, mux_in_sin190, mux_in_cos191, mux_in_sin191, mux_in_cos192, mux_in_sin192, mux_in_cos193, mux_in_sin193, mux_in_cos194, mux_in_sin194, mux_in_cos195, mux_in_sin195, mux_in_cos196, mux_in_sin196, mux_in_cos197, mux_in_sin197, mux_in_cos198, mux_in_sin198, mux_in_cos199, mux_in_sin199, mux_in_cos200, mux_in_sin200, mux_in_cos201, mux_in_sin201, mux_in_cos202, mux_in_sin202, mux_in_cos203, mux_in_sin203, mux_in_cos204, mux_in_sin204, mux_in_cos205, mux_in_sin205, mux_in_cos206, mux_in_sin206, mux_in_cos207, mux_in_sin207, mux_in_cos208, mux_in_sin208, mux_in_cos209, mux_in_sin209, mux_in_cos210, mux_in_sin210, mux_in_cos211, mux_in_sin211, mux_in_cos212, mux_in_sin212, mux_in_cos213, mux_in_sin213, mux_in_cos214, mux_in_sin214, mux_in_cos215, mux_in_sin215, mux_in_cos216, mux_in_sin216, mux_in_cos217, mux_in_sin217, mux_in_cos218, mux_in_sin218, mux_in_cos219, mux_in_sin219, mux_in_cos220, mux_in_sin220, mux_in_cos221, mux_in_sin221, mux_in_cos222, mux_in_sin222, mux_in_cos223, mux_in_sin223, mux_in_cos224, mux_in_sin224, mux_in_cos225, mux_in_sin225, mux_in_cos226, mux_in_sin226, mux_in_cos227, mux_in_sin227, mux_in_cos228, mux_in_sin228, mux_in_cos229, mux_in_sin229, mux_in_cos230, mux_in_sin230, mux_in_cos231, mux_in_sin231, mux_in_cos232, mux_in_sin232, mux_in_cos233, mux_in_sin233, mux_in_cos234, mux_in_sin234, mux_in_cos235, mux_in_sin235, mux_in_cos236, mux_in_sin236, mux_in_cos237, mux_in_sin237, mux_in_cos238, mux_in_sin238, mux_in_cos239, mux_in_sin239, mux_in_cos240, mux_in_sin240, mux_in_cos241, mux_in_sin241, mux_in_cos242, mux_in_sin242, mux_in_cos243, mux_in_sin243, mux_in_cos244, mux_in_sin244, mux_in_cos245, mux_in_sin245, mux_in_cos246, mux_in_sin246, mux_in_cos247, mux_in_sin247, mux_in_cos248, mux_in_sin248, mux_in_cos249, mux_in_sin249, mux_in_cos250, mux_in_sin250, mux_in_cos251, mux_in_sin251, mux_in_cos252, mux_in_sin252, mux_in_cos253, mux_in_sin253, mux_in_cos254, mux_in_sin254, mux_in_cos255, mux_in_sin255, mux_in_cos256, mux_in_sin256, mux_in_cos257, mux_in_sin257, mux_in_cos258, mux_in_sin258, mux_in_cos259, mux_in_sin259, mux_in_cos260, mux_in_sin260, mux_in_cos261, mux_in_sin261, mux_in_cos262, mux_in_sin262, mux_in_cos263, mux_in_sin263, mux_in_cos264, mux_in_sin264, mux_in_cos265, mux_in_sin265, mux_in_cos266, mux_in_sin266, mux_in_cos267, mux_in_sin267, mux_in_cos268, mux_in_sin268, mux_in_cos269, mux_in_sin269, mux_in_cos270, mux_in_sin270, mux_in_cos271, mux_in_sin271, mux_in_cos272, mux_in_sin272, mux_in_cos273, mux_in_sin273, mux_in_cos274, mux_in_sin274, mux_in_cos275, mux_in_sin275, mux_in_cos276, mux_in_sin276, mux_in_cos277, mux_in_sin277, mux_in_cos278, mux_in_sin278, mux_in_cos279, mux_in_sin279, mux_in_cos280, mux_in_sin280, mux_in_cos281, mux_in_sin281, mux_in_cos282, mux_in_sin282, mux_in_cos283, mux_in_sin283, mux_in_cos284, mux_in_sin284, mux_in_cos285, mux_in_sin285, mux_in_cos286, mux_in_sin286, mux_in_cos287, mux_in_sin287, mux_in_cos288, mux_in_sin288, mux_in_cos289, mux_in_sin289, mux_in_cos290, mux_in_sin290, mux_in_cos291, mux_in_sin291, mux_in_cos292, mux_in_sin292, mux_in_cos293, mux_in_sin293, mux_in_cos294, mux_in_sin294, mux_in_cos295, mux_in_sin295, mux_in_cos296, mux_in_sin296, mux_in_cos297, mux_in_sin297, mux_in_cos298, mux_in_sin298, mux_in_cos299, mux_in_sin299, mux_in_cos300, mux_in_sin300, mux_in_cos301, mux_in_sin301, mux_in_cos302, mux_in_sin302, mux_in_cos303, mux_in_sin303, mux_in_cos304, mux_in_sin304, mux_in_cos305, mux_in_sin305, mux_in_cos306, mux_in_sin306, mux_in_cos307, mux_in_sin307, mux_in_cos308, mux_in_sin308, mux_in_cos309, mux_in_sin309, mux_in_cos310, mux_in_sin310, mux_in_cos311, mux_in_sin311, mux_in_cos312, mux_in_sin312, mux_in_cos313, mux_in_sin313, mux_in_cos314, mux_in_sin314, mux_in_cos315, mux_in_sin315, mux_in_cos316, mux_in_sin316, mux_in_cos317, mux_in_sin317, mux_in_cos318, mux_in_sin318, mux_in_cos319, mux_in_sin319, mux_in_cos320, mux_in_sin320, mux_in_cos321, mux_in_sin321, mux_in_cos322, mux_in_sin322, mux_in_cos323, mux_in_sin323, mux_in_cos324, mux_in_sin324, mux_in_cos325, mux_in_sin325, mux_in_cos326, mux_in_sin326, mux_in_cos327, mux_in_sin327, mux_in_cos328, mux_in_sin328, mux_in_cos329, mux_in_sin329, mux_in_cos330, mux_in_sin330, mux_in_cos331, mux_in_sin331, mux_in_cos332, mux_in_sin332, mux_in_cos333, mux_in_sin333, mux_in_cos334, mux_in_sin334, mux_in_cos335, mux_in_sin335, mux_in_cos336, mux_in_sin336, mux_in_cos337, mux_in_sin337, mux_in_cos338, mux_in_sin338, mux_in_cos339, mux_in_sin339, mux_in_cos340, mux_in_sin340, mux_in_cos341, mux_in_sin341, mux_in_cos342, mux_in_sin342, mux_in_cos343, mux_in_sin343, mux_in_cos344, mux_in_sin344, mux_in_cos345, mux_in_sin345, mux_in_cos346, mux_in_sin346, mux_in_cos347, mux_in_sin347, mux_in_cos348, mux_in_sin348, mux_in_cos349, mux_in_sin349, mux_in_cos350, mux_in_sin350, mux_in_cos351, mux_in_sin351, mux_in_cos352, mux_in_sin352, mux_in_cos353, mux_in_sin353, mux_in_cos354, mux_in_sin354, mux_in_cos355, mux_in_sin355, mux_in_cos356, mux_in_sin356, mux_in_cos357, mux_in_sin357, mux_in_cos358, mux_in_sin358, mux_in_cos359, mux_in_sin359, mux_in_cos360, mux_in_sin360, mux_in_cos361, mux_in_sin361, mux_in_cos362, mux_in_sin362, mux_in_cos363, mux_in_sin363, mux_in_cos364, mux_in_sin364, mux_in_cos365, mux_in_sin365, mux_in_cos366, mux_in_sin366, mux_in_cos367, mux_in_sin367, mux_in_cos368, mux_in_sin368, mux_in_cos369, mux_in_sin369, mux_in_cos370, mux_in_sin370, mux_in_cos371, mux_in_sin371, mux_in_cos372, mux_in_sin372, mux_in_cos373, mux_in_sin373, mux_in_cos374, mux_in_sin374, mux_in_cos375, mux_in_sin375, mux_in_cos376, mux_in_sin376, mux_in_cos377, mux_in_sin377, mux_in_cos378, mux_in_sin378, mux_in_cos379, mux_in_sin379, mux_in_cos380, mux_in_sin380, mux_in_cos381, mux_in_sin381, mux_in_cos382, mux_in_sin382, mux_in_cos383, mux_in_sin383, mux_in_cos384, mux_in_sin384, mux_in_cos385, mux_in_sin385, mux_in_cos386, mux_in_sin386, mux_in_cos387, mux_in_sin387, mux_in_cos388, mux_in_sin388, mux_in_cos389, mux_in_sin389, mux_in_cos390, mux_in_sin390, mux_in_cos391, mux_in_sin391, mux_in_cos392, mux_in_sin392, mux_in_cos393, mux_in_sin393, mux_in_cos394, mux_in_sin394, mux_in_cos395, mux_in_sin395, mux_in_cos396, mux_in_sin396, mux_in_cos397, mux_in_sin397, mux_in_cos398, mux_in_sin398, mux_in_cos399, mux_in_sin399, mux_in_cos400, mux_in_sin400, mux_in_cos401, mux_in_sin401, mux_in_cos402, mux_in_sin402, mux_in_cos403, mux_in_sin403, mux_in_cos404, mux_in_sin404, mux_in_cos405, mux_in_sin405, mux_in_cos406, mux_in_sin406, mux_in_cos407, mux_in_sin407, mux_in_cos408, mux_in_sin408, mux_in_cos409, mux_in_sin409, mux_in_cos410, mux_in_sin410, mux_in_cos411, mux_in_sin411, mux_in_cos412, mux_in_sin412, mux_in_cos413, mux_in_sin413, mux_in_cos414, mux_in_sin414, mux_in_cos415, mux_in_sin415, mux_in_cos416, mux_in_sin416, mux_in_cos417, mux_in_sin417, mux_in_cos418, mux_in_sin418, mux_in_cos419, mux_in_sin419, mux_in_cos420, mux_in_sin420, mux_in_cos421, mux_in_sin421, mux_in_cos422, mux_in_sin422, mux_in_cos423, mux_in_sin423, mux_in_cos424, mux_in_sin424, mux_in_cos425, mux_in_sin425, mux_in_cos426, mux_in_sin426, mux_in_cos427, mux_in_sin427, mux_in_cos428, mux_in_sin428, mux_in_cos429, mux_in_sin429, mux_in_cos430, mux_in_sin430, mux_in_cos431, mux_in_sin431, mux_in_cos432, mux_in_sin432, mux_in_cos433, mux_in_sin433, mux_in_cos434, mux_in_sin434, mux_in_cos435, mux_in_sin435, mux_in_cos436, mux_in_sin436, mux_in_cos437, mux_in_sin437, mux_in_cos438, mux_in_sin438, mux_in_cos439, mux_in_sin439, mux_in_cos440, mux_in_sin440, mux_in_cos441, mux_in_sin441, mux_in_cos442, mux_in_sin442, mux_in_cos443, mux_in_sin443, mux_in_cos444, mux_in_sin444, mux_in_cos445, mux_in_sin445, mux_in_cos446, mux_in_sin446, mux_in_cos447, mux_in_sin447, mux_in_cos448, mux_in_sin448, mux_in_cos449, mux_in_sin449, mux_in_cos450, mux_in_sin450, mux_in_cos451, mux_in_sin451, mux_in_cos452, mux_in_sin452, mux_in_cos453, mux_in_sin453, mux_in_cos454, mux_in_sin454, mux_in_cos455, mux_in_sin455, mux_in_cos456, mux_in_sin456, mux_in_cos457, mux_in_sin457, mux_in_cos458, mux_in_sin458, mux_in_cos459, mux_in_sin459, mux_in_cos460, mux_in_sin460, mux_in_cos461, mux_in_sin461, mux_in_cos462, mux_in_sin462, mux_in_cos463, mux_in_sin463, mux_in_cos464, mux_in_sin464, mux_in_cos465, mux_in_sin465, mux_in_cos466, mux_in_sin466, mux_in_cos467, mux_in_sin467, mux_in_cos468, mux_in_sin468, mux_in_cos469, mux_in_sin469, mux_in_cos470, mux_in_sin470, mux_in_cos471, mux_in_sin471, mux_in_cos472, mux_in_sin472, mux_in_cos473, mux_in_sin473, mux_in_cos474, mux_in_sin474, mux_in_cos475, mux_in_sin475, mux_in_cos476, mux_in_sin476, mux_in_cos477, mux_in_sin477, mux_in_cos478, mux_in_sin478, mux_in_cos479, mux_in_sin479, mux_in_cos480, mux_in_sin480, mux_in_cos481, mux_in_sin481, mux_in_cos482, mux_in_sin482, mux_in_cos483, mux_in_sin483, mux_in_cos484, mux_in_sin484, mux_in_cos485, mux_in_sin485, mux_in_cos486, mux_in_sin486, mux_in_cos487, mux_in_sin487, mux_in_cos488, mux_in_sin488, mux_in_cos489, mux_in_sin489, mux_in_cos490, mux_in_sin490, mux_in_cos491, mux_in_sin491, mux_in_cos492, mux_in_sin492, mux_in_cos493, mux_in_sin493, mux_in_cos494, mux_in_sin494, mux_in_cos495, mux_in_sin495, mux_in_cos496, mux_in_sin496, mux_in_cos497, mux_in_sin497, mux_in_cos498, mux_in_sin498, mux_in_cos499, mux_in_sin499, mux_in_cos500, mux_in_sin500, mux_in_cos501, mux_in_sin501, mux_in_cos502, mux_in_sin502, mux_in_cos503, mux_in_sin503, mux_in_cos504, mux_in_sin504, mux_in_cos505, mux_in_sin505, mux_in_cos506, mux_in_sin506, mux_in_cos507, mux_in_sin507, mux_in_cos508, mux_in_sin508, mux_in_cos509, mux_in_sin509, mux_in_cos510, mux_in_sin510, mux_in_cos511, mux_in_sin511, mux_in_cos512, mux_in_sin512;

    assign mux_in_cos0 = 16'b0000000000000000;
    assign mux_in_sin0 = 16'b0000000000000000;
    assign mux_in_cos1 = 16'b0000000000000000;
    assign mux_in_sin1 = 16'b1000000000000000;
    assign mux_in_cos2 = 16'b0000000000000000;
    assign mux_in_sin2 = 16'b1000101001101100;
    assign mux_in_cos3 = 16'b0000000000000000;
    assign mux_in_sin3 = 16'b1001001111001000;
    assign mux_in_cos4 = 16'b0000000000000000;
    assign mux_in_sin4 = 16'b1001101001101100;
    assign mux_in_cos5 = 16'b1111111111111111;
    assign mux_in_sin5 = 16'b1001111110010011;
    assign mux_in_cos6 = 16'b1111111111111111;
    assign mux_in_sin6 = 16'b1010001111001000;
    assign mux_in_cos7 = 16'b1111111111111111;
    assign mux_in_sin7 = 16'b1010011101010111;
    assign mux_in_cos8 = 16'b1111111111111110;
    assign mux_in_sin8 = 16'b1010101001101100;
    assign mux_in_cos9 = 16'b1111111111111110;
    assign mux_in_sin9 = 16'b1010110100100100;
    assign mux_in_cos10 = 16'b1111111111111101;
    assign mux_in_sin10 = 16'b1010111110010010;
    assign mux_in_cos11 = 16'b1111111111111101;
    assign mux_in_sin11 = 16'b1011000111000101;
    assign mux_in_cos12 = 16'b1111111111111100;
    assign mux_in_sin12 = 16'b1011001111000111;
    assign mux_in_cos13 = 16'b1111111111111011;
    assign mux_in_sin13 = 16'b1011010110100000;
    assign mux_in_cos14 = 16'b1111111111111011;
    assign mux_in_sin14 = 16'b1011011101010110;
    assign mux_in_cos15 = 16'b1111111111111010;
    assign mux_in_sin15 = 16'b1011100011101101;
    assign mux_in_cos16 = 16'b1111111111111001;
    assign mux_in_sin16 = 16'b1011101001101010;
    assign mux_in_cos17 = 16'b1111111111111000;
    assign mux_in_sin17 = 16'b1011101111010000;
    assign mux_in_cos18 = 16'b1111111111110111;
    assign mux_in_sin18 = 16'b1011110100100010;
    assign mux_in_cos19 = 16'b1111111111110110;
    assign mux_in_sin19 = 16'b1011111001100001;
    assign mux_in_cos20 = 16'b1111111111110101;
    assign mux_in_sin20 = 16'b1011111110001111;
    assign mux_in_cos21 = 16'b1111111111110100;
    assign mux_in_sin21 = 16'b1100000010101111;
    assign mux_in_cos22 = 16'b1111111111110011;
    assign mux_in_sin22 = 16'b1100000111000010;
    assign mux_in_cos23 = 16'b1111111111110001;
    assign mux_in_sin23 = 16'b1100001011001000;
    assign mux_in_cos24 = 16'b1111111111110000;
    assign mux_in_sin24 = 16'b1100001111000011;
    assign mux_in_cos25 = 16'b1111111111101111;
    assign mux_in_sin25 = 16'b1100010010110100;
    assign mux_in_cos26 = 16'b1111111111101101;
    assign mux_in_sin26 = 16'b1100010110011011;
    assign mux_in_cos27 = 16'b1111111111101100;
    assign mux_in_sin27 = 16'b1100011001111010;
    assign mux_in_cos28 = 16'b1111111111101010;
    assign mux_in_sin28 = 16'b1100011101010000;
    assign mux_in_cos29 = 16'b1111111111101001;
    assign mux_in_sin29 = 16'b1100100000011111;
    assign mux_in_cos30 = 16'b1111111111100111;
    assign mux_in_sin30 = 16'b1100100011100111;
    assign mux_in_cos31 = 16'b1111111111100101;
    assign mux_in_sin31 = 16'b1100100110101000;
    assign mux_in_cos32 = 16'b1111111111100011;
    assign mux_in_sin32 = 16'b1100101001100011;
    assign mux_in_cos33 = 16'b1111111111100010;
    assign mux_in_sin33 = 16'b1100101100011000;
    assign mux_in_cos34 = 16'b1111111111100000;
    assign mux_in_sin34 = 16'b1100101111001000;
    assign mux_in_cos35 = 16'b1111111111011110;
    assign mux_in_sin35 = 16'b1100110001110011;
    assign mux_in_cos36 = 16'b1111111111011100;
    assign mux_in_sin36 = 16'b1100110100011001;
    assign mux_in_cos37 = 16'b1111111111011010;
    assign mux_in_sin37 = 16'b1100110110111010;
    assign mux_in_cos38 = 16'b1111111111011000;
    assign mux_in_sin38 = 16'b1100111001010111;
    assign mux_in_cos39 = 16'b1111111111010110;
    assign mux_in_sin39 = 16'b1100111011101111;
    assign mux_in_cos40 = 16'b1111111111010011;
    assign mux_in_sin40 = 16'b1100111110000100;
    assign mux_in_cos41 = 16'b1111111111010001;
    assign mux_in_sin41 = 16'b1101000000010101;
    assign mux_in_cos42 = 16'b1111111111001111;
    assign mux_in_sin42 = 16'b1101000010100011;
    assign mux_in_cos43 = 16'b1111111111001100;
    assign mux_in_sin43 = 16'b1101000100101101;
    assign mux_in_cos44 = 16'b1111111111001010;
    assign mux_in_sin44 = 16'b1101000110110100;
    assign mux_in_cos45 = 16'b1111111111001000;
    assign mux_in_sin45 = 16'b1101001000111000;
    assign mux_in_cos46 = 16'b1111111111000101;
    assign mux_in_sin46 = 16'b1101001010111001;
    assign mux_in_cos47 = 16'b1111111111000010;
    assign mux_in_sin47 = 16'b1101001100111000;
    assign mux_in_cos48 = 16'b1111111111000000;
    assign mux_in_sin48 = 16'b1101001110110011;
    assign mux_in_cos49 = 16'b1111111110111101;
    assign mux_in_sin49 = 16'b1101010000101100;
    assign mux_in_cos50 = 16'b1111111110111010;
    assign mux_in_sin50 = 16'b1101010010100011;
    assign mux_in_cos51 = 16'b1111111110110111;
    assign mux_in_sin51 = 16'b1101010100010111;
    assign mux_in_cos52 = 16'b1111111110110100;
    assign mux_in_sin52 = 16'b1101010110001000;
    assign mux_in_cos53 = 16'b1111111110110010;
    assign mux_in_sin53 = 16'b1101010111111000;
    assign mux_in_cos54 = 16'b1111111110101111;
    assign mux_in_sin54 = 16'b1101011001100101;
    assign mux_in_cos55 = 16'b1111111110101011;
    assign mux_in_sin55 = 16'b1101011011010001;
    assign mux_in_cos56 = 16'b1111111110101000;
    assign mux_in_sin56 = 16'b1101011100111010;
    assign mux_in_cos57 = 16'b1111111110100101;
    assign mux_in_sin57 = 16'b1101011110100010;
    assign mux_in_cos58 = 16'b1111111110100010;
    assign mux_in_sin58 = 16'b1101100000001000;
    assign mux_in_cos59 = 16'b1111111110011111;
    assign mux_in_sin59 = 16'b1101100001101100;
    assign mux_in_cos60 = 16'b1111111110011011;
    assign mux_in_sin60 = 16'b1101100011001110;
    assign mux_in_cos61 = 16'b1111111110011000;
    assign mux_in_sin61 = 16'b1101100100101110;
    assign mux_in_cos62 = 16'b1111111110010100;
    assign mux_in_sin62 = 16'b1101100110001101;
    assign mux_in_cos63 = 16'b1111111110010001;
    assign mux_in_sin63 = 16'b1101100111101011;
    assign mux_in_cos64 = 16'b1111111110001101;
    assign mux_in_sin64 = 16'b1101101001000111;
    assign mux_in_cos65 = 16'b1111111110001010;
    assign mux_in_sin65 = 16'b1101101010100001;
    assign mux_in_cos66 = 16'b1111111110000110;
    assign mux_in_sin66 = 16'b1101101011111010;
    assign mux_in_cos67 = 16'b1111111110000010;
    assign mux_in_sin67 = 16'b1101101101010010;
    assign mux_in_cos68 = 16'b1111111101111110;
    assign mux_in_sin68 = 16'b1101101110101000;
    assign mux_in_cos69 = 16'b1111111101111011;
    assign mux_in_sin69 = 16'b1101101111111101;
    assign mux_in_cos70 = 16'b1111111101110111;
    assign mux_in_sin70 = 16'b1101110001010001;
    assign mux_in_cos71 = 16'b1111111101110011;
    assign mux_in_sin71 = 16'b1101110010100011;
    assign mux_in_cos72 = 16'b1111111101101111;
    assign mux_in_sin72 = 16'b1101110011110100;
    assign mux_in_cos73 = 16'b1111111101101011;
    assign mux_in_sin73 = 16'b1101110101000101;
    assign mux_in_cos74 = 16'b1111111101100110;
    assign mux_in_sin74 = 16'b1101110110010100;
    assign mux_in_cos75 = 16'b1111111101100010;
    assign mux_in_sin75 = 16'b1101110111100010;
    assign mux_in_cos76 = 16'b1111111101011110;
    assign mux_in_sin76 = 16'b1101111000101110;
    assign mux_in_cos77 = 16'b1111111101011010;
    assign mux_in_sin77 = 16'b1101111001111010;
    assign mux_in_cos78 = 16'b1111111101010101;
    assign mux_in_sin78 = 16'b1101111011000101;
    assign mux_in_cos79 = 16'b1111111101010001;
    assign mux_in_sin79 = 16'b1101111100001111;
    assign mux_in_cos80 = 16'b1111111101001100;
    assign mux_in_sin80 = 16'b1101111101011000;
    assign mux_in_cos81 = 16'b1111111101001000;
    assign mux_in_sin81 = 16'b1101111110100000;
    assign mux_in_cos82 = 16'b1111111101000011;
    assign mux_in_sin82 = 16'b1101111111100111;
    assign mux_in_cos83 = 16'b1111111100111110;
    assign mux_in_sin83 = 16'b1110000000101101;
    assign mux_in_cos84 = 16'b1111111100111010;
    assign mux_in_sin84 = 16'b1110000001110010;
    assign mux_in_cos85 = 16'b1111111100110101;
    assign mux_in_sin85 = 16'b1110000010110110;
    assign mux_in_cos86 = 16'b1111111100110000;
    assign mux_in_sin86 = 16'b1110000011111010;
    assign mux_in_cos87 = 16'b1111111100101011;
    assign mux_in_sin87 = 16'b1110000100111100;
    assign mux_in_cos88 = 16'b1111111100100110;
    assign mux_in_sin88 = 16'b1110000101111110;
    assign mux_in_cos89 = 16'b1111111100100001;
    assign mux_in_sin89 = 16'b1110000111000000;
    assign mux_in_cos90 = 16'b1111111100011100;
    assign mux_in_sin90 = 16'b1110001000000000;
    assign mux_in_cos91 = 16'b1111111100010111;
    assign mux_in_sin91 = 16'b1110001000111111;
    assign mux_in_cos92 = 16'b1111111100010001;
    assign mux_in_sin92 = 16'b1110001001111110;
    assign mux_in_cos93 = 16'b1111111100001100;
    assign mux_in_sin93 = 16'b1110001010111101;
    assign mux_in_cos94 = 16'b1111111100000111;
    assign mux_in_sin94 = 16'b1110001011111010;
    assign mux_in_cos95 = 16'b1111111100000001;
    assign mux_in_sin95 = 16'b1110001100110111;
    assign mux_in_cos96 = 16'b1111111011111100;
    assign mux_in_sin96 = 16'b1110001101110011;
    assign mux_in_cos97 = 16'b1111111011110110;
    assign mux_in_sin97 = 16'b1110001110101110;
    assign mux_in_cos98 = 16'b1111111011110001;
    assign mux_in_sin98 = 16'b1110001111101001;
    assign mux_in_cos99 = 16'b1111111011101011;
    assign mux_in_sin99 = 16'b1110010000100011;
    assign mux_in_cos100 = 16'b1111111011100101;
    assign mux_in_sin100 = 16'b1110010001011101;
    assign mux_in_cos101 = 16'b1111111011100000;
    assign mux_in_sin101 = 16'b1110010010010110;
    assign mux_in_cos102 = 16'b1111111011011010;
    assign mux_in_sin102 = 16'b1110010011001110;
    assign mux_in_cos103 = 16'b1111111011010100;
    assign mux_in_sin103 = 16'b1110010100000110;
    assign mux_in_cos104 = 16'b1111111011001110;
    assign mux_in_sin104 = 16'b1110010100111101;
    assign mux_in_cos105 = 16'b1111111011001000;
    assign mux_in_sin105 = 16'b1110010101110100;
    assign mux_in_cos106 = 16'b1111111011000010;
    assign mux_in_sin106 = 16'b1110010110101010;
    assign mux_in_cos107 = 16'b1111111010111100;
    assign mux_in_sin107 = 16'b1110010111011111;
    assign mux_in_cos108 = 16'b1111111010110110;
    assign mux_in_sin108 = 16'b1110011000010100;
    assign mux_in_cos109 = 16'b1111111010101111;
    assign mux_in_sin109 = 16'b1110011001001000;
    assign mux_in_cos110 = 16'b1111111010101001;
    assign mux_in_sin110 = 16'b1110011001111100;
    assign mux_in_cos111 = 16'b1111111010100011;
    assign mux_in_sin111 = 16'b1110011010110000;
    assign mux_in_cos112 = 16'b1111111010011100;
    assign mux_in_sin112 = 16'b1110011011100011;
    assign mux_in_cos113 = 16'b1111111010010110;
    assign mux_in_sin113 = 16'b1110011100010101;
    assign mux_in_cos114 = 16'b1111111010001111;
    assign mux_in_sin114 = 16'b1110011101000111;
    assign mux_in_cos115 = 16'b1111111010001000;
    assign mux_in_sin115 = 16'b1110011101111001;
    assign mux_in_cos116 = 16'b1111111010000010;
    assign mux_in_sin116 = 16'b1110011110101010;
    assign mux_in_cos117 = 16'b1111111001111011;
    assign mux_in_sin117 = 16'b1110011111011010;
    assign mux_in_cos118 = 16'b1111111001110100;
    assign mux_in_sin118 = 16'b1110100000001010;
    assign mux_in_cos119 = 16'b1111111001101101;
    assign mux_in_sin119 = 16'b1110100000111010;
    assign mux_in_cos120 = 16'b1111111001100110;
    assign mux_in_sin120 = 16'b1110100001101001;
    assign mux_in_cos121 = 16'b1111111001011111;
    assign mux_in_sin121 = 16'b1110100010011000;
    assign mux_in_cos122 = 16'b1111111001011000;
    assign mux_in_sin122 = 16'b1110100011000110;
    assign mux_in_cos123 = 16'b1111111001010001;
    assign mux_in_sin123 = 16'b1110100011110100;
    assign mux_in_cos124 = 16'b1111111001001010;
    assign mux_in_sin124 = 16'b1110100100100010;
    assign mux_in_cos125 = 16'b1111111001000010;
    assign mux_in_sin125 = 16'b1110100101001111;
    assign mux_in_cos126 = 16'b1111111000111011;
    assign mux_in_sin126 = 16'b1110100101111100;
    assign mux_in_cos127 = 16'b1111111000110100;
    assign mux_in_sin127 = 16'b1110100110101000;
    assign mux_in_cos128 = 16'b1111111000101100;
    assign mux_in_sin128 = 16'b1110100111010100;
    assign mux_in_cos129 = 16'b1111111000100101;
    assign mux_in_sin129 = 16'b1110100111111111;
    assign mux_in_cos130 = 16'b1111111000011101;
    assign mux_in_sin130 = 16'b1110101000101011;
    assign mux_in_cos131 = 16'b1111111000010101;
    assign mux_in_sin131 = 16'b1110101001010101;
    assign mux_in_cos132 = 16'b1111111000001110;
    assign mux_in_sin132 = 16'b1110101010000000;
    assign mux_in_cos133 = 16'b1111111000000110;
    assign mux_in_sin133 = 16'b1110101010101010;
    assign mux_in_cos134 = 16'b1111110111111110;
    assign mux_in_sin134 = 16'b1110101011010100;
    assign mux_in_cos135 = 16'b1111110111110110;
    assign mux_in_sin135 = 16'b1110101011111101;
    assign mux_in_cos136 = 16'b1111110111101110;
    assign mux_in_sin136 = 16'b1110101100100110;
    assign mux_in_cos137 = 16'b1111110111100110;
    assign mux_in_sin137 = 16'b1110101101001111;
    assign mux_in_cos138 = 16'b1111110111011110;
    assign mux_in_sin138 = 16'b1110101101110111;
    assign mux_in_cos139 = 16'b1111110111010110;
    assign mux_in_sin139 = 16'b1110101110100000;
    assign mux_in_cos140 = 16'b1111110111001101;
    assign mux_in_sin140 = 16'b1110101111000111;
    assign mux_in_cos141 = 16'b1111110111000101;
    assign mux_in_sin141 = 16'b1110101111101111;
    assign mux_in_cos142 = 16'b1111110110111101;
    assign mux_in_sin142 = 16'b1110110000010110;
    assign mux_in_cos143 = 16'b1111110110110100;
    assign mux_in_sin143 = 16'b1110110000111101;
    assign mux_in_cos144 = 16'b1111110110101100;
    assign mux_in_sin144 = 16'b1110110001100011;
    assign mux_in_cos145 = 16'b1111110110100011;
    assign mux_in_sin145 = 16'b1110110010001001;
    assign mux_in_cos146 = 16'b1111110110011010;
    assign mux_in_sin146 = 16'b1110110010101111;
    assign mux_in_cos147 = 16'b1111110110010001;
    assign mux_in_sin147 = 16'b1110110011010101;
    assign mux_in_cos148 = 16'b1111110110001001;
    assign mux_in_sin148 = 16'b1110110011111010;
    assign mux_in_cos149 = 16'b1111110110000000;
    assign mux_in_sin149 = 16'b1110110100011111;
    assign mux_in_cos150 = 16'b1111110101110111;
    assign mux_in_sin150 = 16'b1110110101000100;
    assign mux_in_cos151 = 16'b1111110101101110;
    assign mux_in_sin151 = 16'b1110110101101000;
    assign mux_in_cos152 = 16'b1111110101100101;
    assign mux_in_sin152 = 16'b1110110110001100;
    assign mux_in_cos153 = 16'b1111110101011100;
    assign mux_in_sin153 = 16'b1110110110110000;
    assign mux_in_cos154 = 16'b1111110101010010;
    assign mux_in_sin154 = 16'b1110110111010100;
    assign mux_in_cos155 = 16'b1111110101001001;
    assign mux_in_sin155 = 16'b1110110111110111;
    assign mux_in_cos156 = 16'b1111110101000000;
    assign mux_in_sin156 = 16'b1110111000011010;
    assign mux_in_cos157 = 16'b1111110100110110;
    assign mux_in_sin157 = 16'b1110111000111101;
    assign mux_in_cos158 = 16'b1111110100101101;
    assign mux_in_sin158 = 16'b1110111001100000;
    assign mux_in_cos159 = 16'b1111110100100011;
    assign mux_in_sin159 = 16'b1110111010000010;
    assign mux_in_cos160 = 16'b1111110100011001;
    assign mux_in_sin160 = 16'b1110111010100100;
    assign mux_in_cos161 = 16'b1111110100010000;
    assign mux_in_sin161 = 16'b1110111011000110;
    assign mux_in_cos162 = 16'b1111110100000110;
    assign mux_in_sin162 = 16'b1110111011100111;
    assign mux_in_cos163 = 16'b1111110011111100;
    assign mux_in_sin163 = 16'b1110111100001001;
    assign mux_in_cos164 = 16'b1111110011110010;
    assign mux_in_sin164 = 16'b1110111100101010;
    assign mux_in_cos165 = 16'b1111110011101000;
    assign mux_in_sin165 = 16'b1110111101001010;
    assign mux_in_cos166 = 16'b1111110011011110;
    assign mux_in_sin166 = 16'b1110111101101011;
    assign mux_in_cos167 = 16'b1111110011010100;
    assign mux_in_sin167 = 16'b1110111110001011;
    assign mux_in_cos168 = 16'b1111110011001010;
    assign mux_in_sin168 = 16'b1110111110101011;
    assign mux_in_cos169 = 16'b1111110010111111;
    assign mux_in_sin169 = 16'b1110111111001011;
    assign mux_in_cos170 = 16'b1111110010110101;
    assign mux_in_sin170 = 16'b1110111111101011;
    assign mux_in_cos171 = 16'b1111110010101011;
    assign mux_in_sin171 = 16'b1111000000001010;
    assign mux_in_cos172 = 16'b1111110010100000;
    assign mux_in_sin172 = 16'b1111000000101010;
    assign mux_in_cos173 = 16'b1111110010010101;
    assign mux_in_sin173 = 16'b1111000001001001;
    assign mux_in_cos174 = 16'b1111110010001011;
    assign mux_in_sin174 = 16'b1111000001100111;
    assign mux_in_cos175 = 16'b1111110010000000;
    assign mux_in_sin175 = 16'b1111000010000110;
    assign mux_in_cos176 = 16'b1111110001110101;
    assign mux_in_sin176 = 16'b1111000010100100;
    assign mux_in_cos177 = 16'b1111110001101010;
    assign mux_in_sin177 = 16'b1111000011000011;
    assign mux_in_cos178 = 16'b1111110001011111;
    assign mux_in_sin178 = 16'b1111000011100000;
    assign mux_in_cos179 = 16'b1111110001010100;
    assign mux_in_sin179 = 16'b1111000011111110;
    assign mux_in_cos180 = 16'b1111110001001001;
    assign mux_in_sin180 = 16'b1111000100011100;
    assign mux_in_cos181 = 16'b1111110000111110;
    assign mux_in_sin181 = 16'b1111000100111001;
    assign mux_in_cos182 = 16'b1111110000110011;
    assign mux_in_sin182 = 16'b1111000101010110;
    assign mux_in_cos183 = 16'b1111110000100111;
    assign mux_in_sin183 = 16'b1111000101110011;
    assign mux_in_cos184 = 16'b1111110000011100;
    assign mux_in_sin184 = 16'b1111000110010000;
    assign mux_in_cos185 = 16'b1111110000010000;
    assign mux_in_sin185 = 16'b1111000110101100;
    assign mux_in_cos186 = 16'b1111110000000101;
    assign mux_in_sin186 = 16'b1111000111001001;
    assign mux_in_cos187 = 16'b1111101111111001;
    assign mux_in_sin187 = 16'b1111000111100101;
    assign mux_in_cos188 = 16'b1111101111101101;
    assign mux_in_sin188 = 16'b1111001000000001;
    assign mux_in_cos189 = 16'b1111101111100001;
    assign mux_in_sin189 = 16'b1111001000011101;
    assign mux_in_cos190 = 16'b1111101111010101;
    assign mux_in_sin190 = 16'b1111001000111000;
    assign mux_in_cos191 = 16'b1111101111001001;
    assign mux_in_sin191 = 16'b1111001001010100;
    assign mux_in_cos192 = 16'b1111101110111101;
    assign mux_in_sin192 = 16'b1111001001101111;
    assign mux_in_cos193 = 16'b1111101110110001;
    assign mux_in_sin193 = 16'b1111001010001010;
    assign mux_in_cos194 = 16'b1111101110100101;
    assign mux_in_sin194 = 16'b1111001010100101;
    assign mux_in_cos195 = 16'b1111101110011001;
    assign mux_in_sin195 = 16'b1111001010111111;
    assign mux_in_cos196 = 16'b1111101110001100;
    assign mux_in_sin196 = 16'b1111001011011010;
    assign mux_in_cos197 = 16'b1111101110000000;
    assign mux_in_sin197 = 16'b1111001011110100;
    assign mux_in_cos198 = 16'b1111101101110011;
    assign mux_in_sin198 = 16'b1111001100001110;
    assign mux_in_cos199 = 16'b1111101101100111;
    assign mux_in_sin199 = 16'b1111001100101000;
    assign mux_in_cos200 = 16'b1111101101011010;
    assign mux_in_sin200 = 16'b1111001101000010;
    assign mux_in_cos201 = 16'b1111101101001101;
    assign mux_in_sin201 = 16'b1111001101011100;
    assign mux_in_cos202 = 16'b1111101101000000;
    assign mux_in_sin202 = 16'b1111001101110101;
    assign mux_in_cos203 = 16'b1111101100110011;
    assign mux_in_sin203 = 16'b1111001110001111;
    assign mux_in_cos204 = 16'b1111101100100110;
    assign mux_in_sin204 = 16'b1111001110101000;
    assign mux_in_cos205 = 16'b1111101100011001;
    assign mux_in_sin205 = 16'b1111001111000001;
    assign mux_in_cos206 = 16'b1111101100001100;
    assign mux_in_sin206 = 16'b1111001111011010;
    assign mux_in_cos207 = 16'b1111101011111110;
    assign mux_in_sin207 = 16'b1111001111110010;
    assign mux_in_cos208 = 16'b1111101011110001;
    assign mux_in_sin208 = 16'b1111010000001011;
    assign mux_in_cos209 = 16'b1111101011100100;
    assign mux_in_sin209 = 16'b1111010000100011;
    assign mux_in_cos210 = 16'b1111101011010110;
    assign mux_in_sin210 = 16'b1111010000111011;
    assign mux_in_cos211 = 16'b1111101011001000;
    assign mux_in_sin211 = 16'b1111010001010100;
    assign mux_in_cos212 = 16'b1111101010111011;
    assign mux_in_sin212 = 16'b1111010001101011;
    assign mux_in_cos213 = 16'b1111101010101101;
    assign mux_in_sin213 = 16'b1111010010000011;
    assign mux_in_cos214 = 16'b1111101010011111;
    assign mux_in_sin214 = 16'b1111010010011011;
    assign mux_in_cos215 = 16'b1111101010010001;
    assign mux_in_sin215 = 16'b1111010010110010;
    assign mux_in_cos216 = 16'b1111101010000011;
    assign mux_in_sin216 = 16'b1111010011001010;
    assign mux_in_cos217 = 16'b1111101001110100;
    assign mux_in_sin217 = 16'b1111010011100001;
    assign mux_in_cos218 = 16'b1111101001100110;
    assign mux_in_sin218 = 16'b1111010011111000;
    assign mux_in_cos219 = 16'b1111101001011000;
    assign mux_in_sin219 = 16'b1111010100001111;
    assign mux_in_cos220 = 16'b1111101001001001;
    assign mux_in_sin220 = 16'b1111010100100101;
    assign mux_in_cos221 = 16'b1111101000111011;
    assign mux_in_sin221 = 16'b1111010100111100;
    assign mux_in_cos222 = 16'b1111101000101100;
    assign mux_in_sin222 = 16'b1111010101010010;
    assign mux_in_cos223 = 16'b1111101000011101;
    assign mux_in_sin223 = 16'b1111010101101001;
    assign mux_in_cos224 = 16'b1111101000001111;
    assign mux_in_sin224 = 16'b1111010101111111;
    assign mux_in_cos225 = 16'b1111101000000000;
    assign mux_in_sin225 = 16'b1111010110010101;
    assign mux_in_cos226 = 16'b1111100111110001;
    assign mux_in_sin226 = 16'b1111010110101011;
    assign mux_in_cos227 = 16'b1111100111100010;
    assign mux_in_sin227 = 16'b1111010111000000;
    assign mux_in_cos228 = 16'b1111100111010010;
    assign mux_in_sin228 = 16'b1111010111010110;
    assign mux_in_cos229 = 16'b1111100111000011;
    assign mux_in_sin229 = 16'b1111010111101100;
    assign mux_in_cos230 = 16'b1111100110110100;
    assign mux_in_sin230 = 16'b1111011000000001;
    assign mux_in_cos231 = 16'b1111100110100100;
    assign mux_in_sin231 = 16'b1111011000010110;
    assign mux_in_cos232 = 16'b1111100110010101;
    assign mux_in_sin232 = 16'b1111011000101011;
    assign mux_in_cos233 = 16'b1111100110000101;
    assign mux_in_sin233 = 16'b1111011001000000;
    assign mux_in_cos234 = 16'b1111100101110101;
    assign mux_in_sin234 = 16'b1111011001010101;
    assign mux_in_cos235 = 16'b1111100101100101;
    assign mux_in_sin235 = 16'b1111011001101010;
    assign mux_in_cos236 = 16'b1111100101010101;
    assign mux_in_sin236 = 16'b1111011001111110;
    assign mux_in_cos237 = 16'b1111100101000101;
    assign mux_in_sin237 = 16'b1111011010010011;
    assign mux_in_cos238 = 16'b1111100100110101;
    assign mux_in_sin238 = 16'b1111011010100111;
    assign mux_in_cos239 = 16'b1111100100100101;
    assign mux_in_sin239 = 16'b1111011010111011;
    assign mux_in_cos240 = 16'b1111100100010100;
    assign mux_in_sin240 = 16'b1111011011001111;
    assign mux_in_cos241 = 16'b1111100100000100;
    assign mux_in_sin241 = 16'b1111011011100011;
    assign mux_in_cos242 = 16'b1111100011110011;
    assign mux_in_sin242 = 16'b1111011011110111;
    assign mux_in_cos243 = 16'b1111100011100011;
    assign mux_in_sin243 = 16'b1111011100001011;
    assign mux_in_cos244 = 16'b1111100011010010;
    assign mux_in_sin244 = 16'b1111011100011110;
    assign mux_in_cos245 = 16'b1111100011000001;
    assign mux_in_sin245 = 16'b1111011100110010;
    assign mux_in_cos246 = 16'b1111100010110000;
    assign mux_in_sin246 = 16'b1111011101000101;
    assign mux_in_cos247 = 16'b1111100010011111;
    assign mux_in_sin247 = 16'b1111011101011000;
    assign mux_in_cos248 = 16'b1111100010001110;
    assign mux_in_sin248 = 16'b1111011101101011;
    assign mux_in_cos249 = 16'b1111100001111100;
    assign mux_in_sin249 = 16'b1111011101111110;
    assign mux_in_cos250 = 16'b1111100001101011;
    assign mux_in_sin250 = 16'b1111011110010001;
    assign mux_in_cos251 = 16'b1111100001011001;
    assign mux_in_sin251 = 16'b1111011110100100;
    assign mux_in_cos252 = 16'b1111100001001000;
    assign mux_in_sin252 = 16'b1111011110110111;
    assign mux_in_cos253 = 16'b1111100000110110;
    assign mux_in_sin253 = 16'b1111011111001001;
    assign mux_in_cos254 = 16'b1111100000100100;
    assign mux_in_sin254 = 16'b1111011111011100;
    assign mux_in_cos255 = 16'b1111100000010010;
    assign mux_in_sin255 = 16'b1111011111101110;
    assign mux_in_cos256 = 16'b1111100000000000;
    assign mux_in_sin256 = 16'b1111100000000000;
    assign mux_in_cos257 = 16'b1111011111101110;
    assign mux_in_sin257 = 16'b1111100000010010;
    assign mux_in_cos258 = 16'b1111011111011100;
    assign mux_in_sin258 = 16'b1111100000100100;
    assign mux_in_cos259 = 16'b1111011111001001;
    assign mux_in_sin259 = 16'b1111100000110110;
    assign mux_in_cos260 = 16'b1111011110110111;
    assign mux_in_sin260 = 16'b1111100001001000;
    assign mux_in_cos261 = 16'b1111011110100100;
    assign mux_in_sin261 = 16'b1111100001011001;
    assign mux_in_cos262 = 16'b1111011110010001;
    assign mux_in_sin262 = 16'b1111100001101011;
    assign mux_in_cos263 = 16'b1111011101111110;
    assign mux_in_sin263 = 16'b1111100001111100;
    assign mux_in_cos264 = 16'b1111011101101011;
    assign mux_in_sin264 = 16'b1111100010001110;
    assign mux_in_cos265 = 16'b1111011101011000;
    assign mux_in_sin265 = 16'b1111100010011111;
    assign mux_in_cos266 = 16'b1111011101000101;
    assign mux_in_sin266 = 16'b1111100010110000;
    assign mux_in_cos267 = 16'b1111011100110010;
    assign mux_in_sin267 = 16'b1111100011000001;
    assign mux_in_cos268 = 16'b1111011100011110;
    assign mux_in_sin268 = 16'b1111100011010010;
    assign mux_in_cos269 = 16'b1111011100001011;
    assign mux_in_sin269 = 16'b1111100011100011;
    assign mux_in_cos270 = 16'b1111011011110111;
    assign mux_in_sin270 = 16'b1111100011110011;
    assign mux_in_cos271 = 16'b1111011011100011;
    assign mux_in_sin271 = 16'b1111100100000100;
    assign mux_in_cos272 = 16'b1111011011001111;
    assign mux_in_sin272 = 16'b1111100100010100;
    assign mux_in_cos273 = 16'b1111011010111011;
    assign mux_in_sin273 = 16'b1111100100100101;
    assign mux_in_cos274 = 16'b1111011010100111;
    assign mux_in_sin274 = 16'b1111100100110101;
    assign mux_in_cos275 = 16'b1111011010010011;
    assign mux_in_sin275 = 16'b1111100101000101;
    assign mux_in_cos276 = 16'b1111011001111110;
    assign mux_in_sin276 = 16'b1111100101010101;
    assign mux_in_cos277 = 16'b1111011001101010;
    assign mux_in_sin277 = 16'b1111100101100101;
    assign mux_in_cos278 = 16'b1111011001010101;
    assign mux_in_sin278 = 16'b1111100101110101;
    assign mux_in_cos279 = 16'b1111011001000000;
    assign mux_in_sin279 = 16'b1111100110000101;
    assign mux_in_cos280 = 16'b1111011000101011;
    assign mux_in_sin280 = 16'b1111100110010101;
    assign mux_in_cos281 = 16'b1111011000010110;
    assign mux_in_sin281 = 16'b1111100110100100;
    assign mux_in_cos282 = 16'b1111011000000001;
    assign mux_in_sin282 = 16'b1111100110110100;
    assign mux_in_cos283 = 16'b1111010111101100;
    assign mux_in_sin283 = 16'b1111100111000011;
    assign mux_in_cos284 = 16'b1111010111010110;
    assign mux_in_sin284 = 16'b1111100111010010;
    assign mux_in_cos285 = 16'b1111010111000000;
    assign mux_in_sin285 = 16'b1111100111100010;
    assign mux_in_cos286 = 16'b1111010110101011;
    assign mux_in_sin286 = 16'b1111100111110001;
    assign mux_in_cos287 = 16'b1111010110010101;
    assign mux_in_sin287 = 16'b1111101000000000;
    assign mux_in_cos288 = 16'b1111010101111111;
    assign mux_in_sin288 = 16'b1111101000001111;
    assign mux_in_cos289 = 16'b1111010101101001;
    assign mux_in_sin289 = 16'b1111101000011101;
    assign mux_in_cos290 = 16'b1111010101010010;
    assign mux_in_sin290 = 16'b1111101000101100;
    assign mux_in_cos291 = 16'b1111010100111100;
    assign mux_in_sin291 = 16'b1111101000111011;
    assign mux_in_cos292 = 16'b1111010100100101;
    assign mux_in_sin292 = 16'b1111101001001001;
    assign mux_in_cos293 = 16'b1111010100001111;
    assign mux_in_sin293 = 16'b1111101001011000;
    assign mux_in_cos294 = 16'b1111010011111000;
    assign mux_in_sin294 = 16'b1111101001100110;
    assign mux_in_cos295 = 16'b1111010011100001;
    assign mux_in_sin295 = 16'b1111101001110100;
    assign mux_in_cos296 = 16'b1111010011001010;
    assign mux_in_sin296 = 16'b1111101010000011;
    assign mux_in_cos297 = 16'b1111010010110010;
    assign mux_in_sin297 = 16'b1111101010010001;
    assign mux_in_cos298 = 16'b1111010010011011;
    assign mux_in_sin298 = 16'b1111101010011111;
    assign mux_in_cos299 = 16'b1111010010000011;
    assign mux_in_sin299 = 16'b1111101010101101;
    assign mux_in_cos300 = 16'b1111010001101011;
    assign mux_in_sin300 = 16'b1111101010111011;
    assign mux_in_cos301 = 16'b1111010001010100;
    assign mux_in_sin301 = 16'b1111101011001000;
    assign mux_in_cos302 = 16'b1111010000111011;
    assign mux_in_sin302 = 16'b1111101011010110;
    assign mux_in_cos303 = 16'b1111010000100011;
    assign mux_in_sin303 = 16'b1111101011100100;
    assign mux_in_cos304 = 16'b1111010000001011;
    assign mux_in_sin304 = 16'b1111101011110001;
    assign mux_in_cos305 = 16'b1111001111110010;
    assign mux_in_sin305 = 16'b1111101011111110;
    assign mux_in_cos306 = 16'b1111001111011010;
    assign mux_in_sin306 = 16'b1111101100001100;
    assign mux_in_cos307 = 16'b1111001111000001;
    assign mux_in_sin307 = 16'b1111101100011001;
    assign mux_in_cos308 = 16'b1111001110101000;
    assign mux_in_sin308 = 16'b1111101100100110;
    assign mux_in_cos309 = 16'b1111001110001111;
    assign mux_in_sin309 = 16'b1111101100110011;
    assign mux_in_cos310 = 16'b1111001101110101;
    assign mux_in_sin310 = 16'b1111101101000000;
    assign mux_in_cos311 = 16'b1111001101011100;
    assign mux_in_sin311 = 16'b1111101101001101;
    assign mux_in_cos312 = 16'b1111001101000010;
    assign mux_in_sin312 = 16'b1111101101011010;
    assign mux_in_cos313 = 16'b1111001100101000;
    assign mux_in_sin313 = 16'b1111101101100111;
    assign mux_in_cos314 = 16'b1111001100001110;
    assign mux_in_sin314 = 16'b1111101101110011;
    assign mux_in_cos315 = 16'b1111001011110100;
    assign mux_in_sin315 = 16'b1111101110000000;
    assign mux_in_cos316 = 16'b1111001011011010;
    assign mux_in_sin316 = 16'b1111101110001100;
    assign mux_in_cos317 = 16'b1111001010111111;
    assign mux_in_sin317 = 16'b1111101110011001;
    assign mux_in_cos318 = 16'b1111001010100101;
    assign mux_in_sin318 = 16'b1111101110100101;
    assign mux_in_cos319 = 16'b1111001010001010;
    assign mux_in_sin319 = 16'b1111101110110001;
    assign mux_in_cos320 = 16'b1111001001101111;
    assign mux_in_sin320 = 16'b1111101110111101;
    assign mux_in_cos321 = 16'b1111001001010100;
    assign mux_in_sin321 = 16'b1111101111001001;
    assign mux_in_cos322 = 16'b1111001000111000;
    assign mux_in_sin322 = 16'b1111101111010101;
    assign mux_in_cos323 = 16'b1111001000011101;
    assign mux_in_sin323 = 16'b1111101111100001;
    assign mux_in_cos324 = 16'b1111001000000001;
    assign mux_in_sin324 = 16'b1111101111101101;
    assign mux_in_cos325 = 16'b1111000111100101;
    assign mux_in_sin325 = 16'b1111101111111001;
    assign mux_in_cos326 = 16'b1111000111001001;
    assign mux_in_sin326 = 16'b1111110000000101;
    assign mux_in_cos327 = 16'b1111000110101100;
    assign mux_in_sin327 = 16'b1111110000010000;
    assign mux_in_cos328 = 16'b1111000110010000;
    assign mux_in_sin328 = 16'b1111110000011100;
    assign mux_in_cos329 = 16'b1111000101110011;
    assign mux_in_sin329 = 16'b1111110000100111;
    assign mux_in_cos330 = 16'b1111000101010110;
    assign mux_in_sin330 = 16'b1111110000110011;
    assign mux_in_cos331 = 16'b1111000100111001;
    assign mux_in_sin331 = 16'b1111110000111110;
    assign mux_in_cos332 = 16'b1111000100011100;
    assign mux_in_sin332 = 16'b1111110001001001;
    assign mux_in_cos333 = 16'b1111000011111110;
    assign mux_in_sin333 = 16'b1111110001010100;
    assign mux_in_cos334 = 16'b1111000011100000;
    assign mux_in_sin334 = 16'b1111110001011111;
    assign mux_in_cos335 = 16'b1111000011000011;
    assign mux_in_sin335 = 16'b1111110001101010;
    assign mux_in_cos336 = 16'b1111000010100100;
    assign mux_in_sin336 = 16'b1111110001110101;
    assign mux_in_cos337 = 16'b1111000010000110;
    assign mux_in_sin337 = 16'b1111110010000000;
    assign mux_in_cos338 = 16'b1111000001100111;
    assign mux_in_sin338 = 16'b1111110010001011;
    assign mux_in_cos339 = 16'b1111000001001001;
    assign mux_in_sin339 = 16'b1111110010010101;
    assign mux_in_cos340 = 16'b1111000000101010;
    assign mux_in_sin340 = 16'b1111110010100000;
    assign mux_in_cos341 = 16'b1111000000001010;
    assign mux_in_sin341 = 16'b1111110010101011;
    assign mux_in_cos342 = 16'b1110111111101011;
    assign mux_in_sin342 = 16'b1111110010110101;
    assign mux_in_cos343 = 16'b1110111111001011;
    assign mux_in_sin343 = 16'b1111110010111111;
    assign mux_in_cos344 = 16'b1110111110101011;
    assign mux_in_sin344 = 16'b1111110011001010;
    assign mux_in_cos345 = 16'b1110111110001011;
    assign mux_in_sin345 = 16'b1111110011010100;
    assign mux_in_cos346 = 16'b1110111101101011;
    assign mux_in_sin346 = 16'b1111110011011110;
    assign mux_in_cos347 = 16'b1110111101001010;
    assign mux_in_sin347 = 16'b1111110011101000;
    assign mux_in_cos348 = 16'b1110111100101010;
    assign mux_in_sin348 = 16'b1111110011110010;
    assign mux_in_cos349 = 16'b1110111100001001;
    assign mux_in_sin349 = 16'b1111110011111100;
    assign mux_in_cos350 = 16'b1110111011100111;
    assign mux_in_sin350 = 16'b1111110100000110;
    assign mux_in_cos351 = 16'b1110111011000110;
    assign mux_in_sin351 = 16'b1111110100010000;
    assign mux_in_cos352 = 16'b1110111010100100;
    assign mux_in_sin352 = 16'b1111110100011001;
    assign mux_in_cos353 = 16'b1110111010000010;
    assign mux_in_sin353 = 16'b1111110100100011;
    assign mux_in_cos354 = 16'b1110111001100000;
    assign mux_in_sin354 = 16'b1111110100101101;
    assign mux_in_cos355 = 16'b1110111000111101;
    assign mux_in_sin355 = 16'b1111110100110110;
    assign mux_in_cos356 = 16'b1110111000011010;
    assign mux_in_sin356 = 16'b1111110101000000;
    assign mux_in_cos357 = 16'b1110110111110111;
    assign mux_in_sin357 = 16'b1111110101001001;
    assign mux_in_cos358 = 16'b1110110111010100;
    assign mux_in_sin358 = 16'b1111110101010010;
    assign mux_in_cos359 = 16'b1110110110110000;
    assign mux_in_sin359 = 16'b1111110101011100;
    assign mux_in_cos360 = 16'b1110110110001100;
    assign mux_in_sin360 = 16'b1111110101100101;
    assign mux_in_cos361 = 16'b1110110101101000;
    assign mux_in_sin361 = 16'b1111110101101110;
    assign mux_in_cos362 = 16'b1110110101000100;
    assign mux_in_sin362 = 16'b1111110101110111;
    assign mux_in_cos363 = 16'b1110110100011111;
    assign mux_in_sin363 = 16'b1111110110000000;
    assign mux_in_cos364 = 16'b1110110011111010;
    assign mux_in_sin364 = 16'b1111110110001001;
    assign mux_in_cos365 = 16'b1110110011010101;
    assign mux_in_sin365 = 16'b1111110110010001;
    assign mux_in_cos366 = 16'b1110110010101111;
    assign mux_in_sin366 = 16'b1111110110011010;
    assign mux_in_cos367 = 16'b1110110010001001;
    assign mux_in_sin367 = 16'b1111110110100011;
    assign mux_in_cos368 = 16'b1110110001100011;
    assign mux_in_sin368 = 16'b1111110110101100;
    assign mux_in_cos369 = 16'b1110110000111101;
    assign mux_in_sin369 = 16'b1111110110110100;
    assign mux_in_cos370 = 16'b1110110000010110;
    assign mux_in_sin370 = 16'b1111110110111101;
    assign mux_in_cos371 = 16'b1110101111101111;
    assign mux_in_sin371 = 16'b1111110111000101;
    assign mux_in_cos372 = 16'b1110101111000111;
    assign mux_in_sin372 = 16'b1111110111001101;
    assign mux_in_cos373 = 16'b1110101110100000;
    assign mux_in_sin373 = 16'b1111110111010110;
    assign mux_in_cos374 = 16'b1110101101110111;
    assign mux_in_sin374 = 16'b1111110111011110;
    assign mux_in_cos375 = 16'b1110101101001111;
    assign mux_in_sin375 = 16'b1111110111100110;
    assign mux_in_cos376 = 16'b1110101100100110;
    assign mux_in_sin376 = 16'b1111110111101110;
    assign mux_in_cos377 = 16'b1110101011111101;
    assign mux_in_sin377 = 16'b1111110111110110;
    assign mux_in_cos378 = 16'b1110101011010100;
    assign mux_in_sin378 = 16'b1111110111111110;
    assign mux_in_cos379 = 16'b1110101010101010;
    assign mux_in_sin379 = 16'b1111111000000110;
    assign mux_in_cos380 = 16'b1110101010000000;
    assign mux_in_sin380 = 16'b1111111000001110;
    assign mux_in_cos381 = 16'b1110101001010101;
    assign mux_in_sin381 = 16'b1111111000010101;
    assign mux_in_cos382 = 16'b1110101000101011;
    assign mux_in_sin382 = 16'b1111111000011101;
    assign mux_in_cos383 = 16'b1110100111111111;
    assign mux_in_sin383 = 16'b1111111000100101;
    assign mux_in_cos384 = 16'b1110100111010100;
    assign mux_in_sin384 = 16'b1111111000101100;
    assign mux_in_cos385 = 16'b1110100110101000;
    assign mux_in_sin385 = 16'b1111111000110100;
    assign mux_in_cos386 = 16'b1110100101111100;
    assign mux_in_sin386 = 16'b1111111000111011;
    assign mux_in_cos387 = 16'b1110100101001111;
    assign mux_in_sin387 = 16'b1111111001000010;
    assign mux_in_cos388 = 16'b1110100100100010;
    assign mux_in_sin388 = 16'b1111111001001010;
    assign mux_in_cos389 = 16'b1110100011110100;
    assign mux_in_sin389 = 16'b1111111001010001;
    assign mux_in_cos390 = 16'b1110100011000110;
    assign mux_in_sin390 = 16'b1111111001011000;
    assign mux_in_cos391 = 16'b1110100010011000;
    assign mux_in_sin391 = 16'b1111111001011111;
    assign mux_in_cos392 = 16'b1110100001101001;
    assign mux_in_sin392 = 16'b1111111001100110;
    assign mux_in_cos393 = 16'b1110100000111010;
    assign mux_in_sin393 = 16'b1111111001101101;
    assign mux_in_cos394 = 16'b1110100000001010;
    assign mux_in_sin394 = 16'b1111111001110100;
    assign mux_in_cos395 = 16'b1110011111011010;
    assign mux_in_sin395 = 16'b1111111001111011;
    assign mux_in_cos396 = 16'b1110011110101010;
    assign mux_in_sin396 = 16'b1111111010000010;
    assign mux_in_cos397 = 16'b1110011101111001;
    assign mux_in_sin397 = 16'b1111111010001000;
    assign mux_in_cos398 = 16'b1110011101000111;
    assign mux_in_sin398 = 16'b1111111010001111;
    assign mux_in_cos399 = 16'b1110011100010101;
    assign mux_in_sin399 = 16'b1111111010010110;
    assign mux_in_cos400 = 16'b1110011011100011;
    assign mux_in_sin400 = 16'b1111111010011100;
    assign mux_in_cos401 = 16'b1110011010110000;
    assign mux_in_sin401 = 16'b1111111010100011;
    assign mux_in_cos402 = 16'b1110011001111100;
    assign mux_in_sin402 = 16'b1111111010101001;
    assign mux_in_cos403 = 16'b1110011001001000;
    assign mux_in_sin403 = 16'b1111111010101111;
    assign mux_in_cos404 = 16'b1110011000010100;
    assign mux_in_sin404 = 16'b1111111010110110;
    assign mux_in_cos405 = 16'b1110010111011111;
    assign mux_in_sin405 = 16'b1111111010111100;
    assign mux_in_cos406 = 16'b1110010110101010;
    assign mux_in_sin406 = 16'b1111111011000010;
    assign mux_in_cos407 = 16'b1110010101110100;
    assign mux_in_sin407 = 16'b1111111011001000;
    assign mux_in_cos408 = 16'b1110010100111101;
    assign mux_in_sin408 = 16'b1111111011001110;
    assign mux_in_cos409 = 16'b1110010100000110;
    assign mux_in_sin409 = 16'b1111111011010100;
    assign mux_in_cos410 = 16'b1110010011001110;
    assign mux_in_sin410 = 16'b1111111011011010;
    assign mux_in_cos411 = 16'b1110010010010110;
    assign mux_in_sin411 = 16'b1111111011100000;
    assign mux_in_cos412 = 16'b1110010001011101;
    assign mux_in_sin412 = 16'b1111111011100101;
    assign mux_in_cos413 = 16'b1110010000100011;
    assign mux_in_sin413 = 16'b1111111011101011;
    assign mux_in_cos414 = 16'b1110001111101001;
    assign mux_in_sin414 = 16'b1111111011110001;
    assign mux_in_cos415 = 16'b1110001110101110;
    assign mux_in_sin415 = 16'b1111111011110110;
    assign mux_in_cos416 = 16'b1110001101110011;
    assign mux_in_sin416 = 16'b1111111011111100;
    assign mux_in_cos417 = 16'b1110001100110111;
    assign mux_in_sin417 = 16'b1111111100000001;
    assign mux_in_cos418 = 16'b1110001011111010;
    assign mux_in_sin418 = 16'b1111111100000111;
    assign mux_in_cos419 = 16'b1110001010111101;
    assign mux_in_sin419 = 16'b1111111100001100;
    assign mux_in_cos420 = 16'b1110001001111110;
    assign mux_in_sin420 = 16'b1111111100010001;
    assign mux_in_cos421 = 16'b1110001000111111;
    assign mux_in_sin421 = 16'b1111111100010111;
    assign mux_in_cos422 = 16'b1110001000000000;
    assign mux_in_sin422 = 16'b1111111100011100;
    assign mux_in_cos423 = 16'b1110000111000000;
    assign mux_in_sin423 = 16'b1111111100100001;
    assign mux_in_cos424 = 16'b1110000101111110;
    assign mux_in_sin424 = 16'b1111111100100110;
    assign mux_in_cos425 = 16'b1110000100111100;
    assign mux_in_sin425 = 16'b1111111100101011;
    assign mux_in_cos426 = 16'b1110000011111010;
    assign mux_in_sin426 = 16'b1111111100110000;
    assign mux_in_cos427 = 16'b1110000010110110;
    assign mux_in_sin427 = 16'b1111111100110101;
    assign mux_in_cos428 = 16'b1110000001110010;
    assign mux_in_sin428 = 16'b1111111100111010;
    assign mux_in_cos429 = 16'b1110000000101101;
    assign mux_in_sin429 = 16'b1111111100111110;
    assign mux_in_cos430 = 16'b1101111111100111;
    assign mux_in_sin430 = 16'b1111111101000011;
    assign mux_in_cos431 = 16'b1101111110100000;
    assign mux_in_sin431 = 16'b1111111101001000;
    assign mux_in_cos432 = 16'b1101111101011000;
    assign mux_in_sin432 = 16'b1111111101001100;
    assign mux_in_cos433 = 16'b1101111100001111;
    assign mux_in_sin433 = 16'b1111111101010001;
    assign mux_in_cos434 = 16'b1101111011000101;
    assign mux_in_sin434 = 16'b1111111101010101;
    assign mux_in_cos435 = 16'b1101111001111010;
    assign mux_in_sin435 = 16'b1111111101011010;
    assign mux_in_cos436 = 16'b1101111000101110;
    assign mux_in_sin436 = 16'b1111111101011110;
    assign mux_in_cos437 = 16'b1101110111100010;
    assign mux_in_sin437 = 16'b1111111101100010;
    assign mux_in_cos438 = 16'b1101110110010100;
    assign mux_in_sin438 = 16'b1111111101100110;
    assign mux_in_cos439 = 16'b1101110101000101;
    assign mux_in_sin439 = 16'b1111111101101011;
    assign mux_in_cos440 = 16'b1101110011110100;
    assign mux_in_sin440 = 16'b1111111101101111;
    assign mux_in_cos441 = 16'b1101110010100011;
    assign mux_in_sin441 = 16'b1111111101110011;
    assign mux_in_cos442 = 16'b1101110001010001;
    assign mux_in_sin442 = 16'b1111111101110111;
    assign mux_in_cos443 = 16'b1101101111111101;
    assign mux_in_sin443 = 16'b1111111101111011;
    assign mux_in_cos444 = 16'b1101101110101000;
    assign mux_in_sin444 = 16'b1111111101111110;
    assign mux_in_cos445 = 16'b1101101101010010;
    assign mux_in_sin445 = 16'b1111111110000010;
    assign mux_in_cos446 = 16'b1101101011111010;
    assign mux_in_sin446 = 16'b1111111110000110;
    assign mux_in_cos447 = 16'b1101101010100001;
    assign mux_in_sin447 = 16'b1111111110001010;
    assign mux_in_cos448 = 16'b1101101001000111;
    assign mux_in_sin448 = 16'b1111111110001101;
    assign mux_in_cos449 = 16'b1101100111101011;
    assign mux_in_sin449 = 16'b1111111110010001;
    assign mux_in_cos450 = 16'b1101100110001101;
    assign mux_in_sin450 = 16'b1111111110010100;
    assign mux_in_cos451 = 16'b1101100100101110;
    assign mux_in_sin451 = 16'b1111111110011000;
    assign mux_in_cos452 = 16'b1101100011001110;
    assign mux_in_sin452 = 16'b1111111110011011;
    assign mux_in_cos453 = 16'b1101100001101100;
    assign mux_in_sin453 = 16'b1111111110011111;
    assign mux_in_cos454 = 16'b1101100000001000;
    assign mux_in_sin454 = 16'b1111111110100010;
    assign mux_in_cos455 = 16'b1101011110100010;
    assign mux_in_sin455 = 16'b1111111110100101;
    assign mux_in_cos456 = 16'b1101011100111010;
    assign mux_in_sin456 = 16'b1111111110101000;
    assign mux_in_cos457 = 16'b1101011011010001;
    assign mux_in_sin457 = 16'b1111111110101011;
    assign mux_in_cos458 = 16'b1101011001100101;
    assign mux_in_sin458 = 16'b1111111110101111;
    assign mux_in_cos459 = 16'b1101010111111000;
    assign mux_in_sin459 = 16'b1111111110110010;
    assign mux_in_cos460 = 16'b1101010110001000;
    assign mux_in_sin460 = 16'b1111111110110100;
    assign mux_in_cos461 = 16'b1101010100010111;
    assign mux_in_sin461 = 16'b1111111110110111;
    assign mux_in_cos462 = 16'b1101010010100011;
    assign mux_in_sin462 = 16'b1111111110111010;
    assign mux_in_cos463 = 16'b1101010000101100;
    assign mux_in_sin463 = 16'b1111111110111101;
    assign mux_in_cos464 = 16'b1101001110110011;
    assign mux_in_sin464 = 16'b1111111111000000;
    assign mux_in_cos465 = 16'b1101001100111000;
    assign mux_in_sin465 = 16'b1111111111000010;
    assign mux_in_cos466 = 16'b1101001010111001;
    assign mux_in_sin466 = 16'b1111111111000101;
    assign mux_in_cos467 = 16'b1101001000111000;
    assign mux_in_sin467 = 16'b1111111111001000;
    assign mux_in_cos468 = 16'b1101000110110100;
    assign mux_in_sin468 = 16'b1111111111001010;
    assign mux_in_cos469 = 16'b1101000100101101;
    assign mux_in_sin469 = 16'b1111111111001100;
    assign mux_in_cos470 = 16'b1101000010100011;
    assign mux_in_sin470 = 16'b1111111111001111;
    assign mux_in_cos471 = 16'b1101000000010101;
    assign mux_in_sin471 = 16'b1111111111010001;
    assign mux_in_cos472 = 16'b1100111110000100;
    assign mux_in_sin472 = 16'b1111111111010011;
    assign mux_in_cos473 = 16'b1100111011101111;
    assign mux_in_sin473 = 16'b1111111111010110;
    assign mux_in_cos474 = 16'b1100111001010111;
    assign mux_in_sin474 = 16'b1111111111011000;
    assign mux_in_cos475 = 16'b1100110110111010;
    assign mux_in_sin475 = 16'b1111111111011010;
    assign mux_in_cos476 = 16'b1100110100011001;
    assign mux_in_sin476 = 16'b1111111111011100;
    assign mux_in_cos477 = 16'b1100110001110011;
    assign mux_in_sin477 = 16'b1111111111011110;
    assign mux_in_cos478 = 16'b1100101111001000;
    assign mux_in_sin478 = 16'b1111111111100000;
    assign mux_in_cos479 = 16'b1100101100011000;
    assign mux_in_sin479 = 16'b1111111111100010;
    assign mux_in_cos480 = 16'b1100101001100011;
    assign mux_in_sin480 = 16'b1111111111100011;
    assign mux_in_cos481 = 16'b1100100110101000;
    assign mux_in_sin481 = 16'b1111111111100101;
    assign mux_in_cos482 = 16'b1100100011100111;
    assign mux_in_sin482 = 16'b1111111111100111;
    assign mux_in_cos483 = 16'b1100100000011111;
    assign mux_in_sin483 = 16'b1111111111101001;
    assign mux_in_cos484 = 16'b1100011101010000;
    assign mux_in_sin484 = 16'b1111111111101010;
    assign mux_in_cos485 = 16'b1100011001111010;
    assign mux_in_sin485 = 16'b1111111111101100;
    assign mux_in_cos486 = 16'b1100010110011011;
    assign mux_in_sin486 = 16'b1111111111101101;
    assign mux_in_cos487 = 16'b1100010010110100;
    assign mux_in_sin487 = 16'b1111111111101111;
    assign mux_in_cos488 = 16'b1100001111000011;
    assign mux_in_sin488 = 16'b1111111111110000;
    assign mux_in_cos489 = 16'b1100001011001000;
    assign mux_in_sin489 = 16'b1111111111110001;
    assign mux_in_cos490 = 16'b1100000111000010;
    assign mux_in_sin490 = 16'b1111111111110011;
    assign mux_in_cos491 = 16'b1100000010101111;
    assign mux_in_sin491 = 16'b1111111111110100;
    assign mux_in_cos492 = 16'b1011111110001111;
    assign mux_in_sin492 = 16'b1111111111110101;
    assign mux_in_cos493 = 16'b1011111001100001;
    assign mux_in_sin493 = 16'b1111111111110110;
    assign mux_in_cos494 = 16'b1011110100100010;
    assign mux_in_sin494 = 16'b1111111111110111;
    assign mux_in_cos495 = 16'b1011101111010000;
    assign mux_in_sin495 = 16'b1111111111111000;
    assign mux_in_cos496 = 16'b1011101001101010;
    assign mux_in_sin496 = 16'b1111111111111001;
    assign mux_in_cos497 = 16'b1011100011101101;
    assign mux_in_sin497 = 16'b1111111111111010;
    assign mux_in_cos498 = 16'b1011011101010110;
    assign mux_in_sin498 = 16'b1111111111111011;
    assign mux_in_cos499 = 16'b1011010110100000;
    assign mux_in_sin499 = 16'b1111111111111011;
    assign mux_in_cos500 = 16'b1011001111000111;
    assign mux_in_sin500 = 16'b1111111111111100;
    assign mux_in_cos501 = 16'b1011000111000101;
    assign mux_in_sin501 = 16'b1111111111111101;
    assign mux_in_cos502 = 16'b1010111110010010;
    assign mux_in_sin502 = 16'b1111111111111101;
    assign mux_in_cos503 = 16'b1010110100100100;
    assign mux_in_sin503 = 16'b1111111111111110;
    assign mux_in_cos504 = 16'b1010101001101100;
    assign mux_in_sin504 = 16'b1111111111111110;
    assign mux_in_cos505 = 16'b1010011101010111;
    assign mux_in_sin505 = 16'b1111111111111111;
    assign mux_in_cos506 = 16'b1010001111001000;
    assign mux_in_sin506 = 16'b1111111111111111;
    assign mux_in_cos507 = 16'b1001111110010011;
    assign mux_in_sin507 = 16'b1111111111111111;
    assign mux_in_cos508 = 16'b1001101001101100;
    assign mux_in_sin508 = 16'b0000000000000000;
    assign mux_in_cos509 = 16'b1001001111001000;
    assign mux_in_sin509 = 16'b0000000000000000;
    assign mux_in_cos510 = 16'b1000101001101100;
    assign mux_in_sin510 = 16'b0000000000000000;
    assign mux_in_cos511 = 16'b1000000000000000;
    assign mux_in_sin511 = 16'b0000000000000000;
    assign mux_in_cos512 = 16'b0000000000000000;
    assign mux_in_sin512 = 16'b0000000000000000;

    always @ (*)
    begin
        case(x_in1)
        10'b0000000000 : logsin1 = mux_in_sin0;
        10'b0000000001 : logsin1 = mux_in_sin1;
        10'b0000000010 : logsin1 = mux_in_sin2;
        10'b0000000011 : logsin1 = mux_in_sin3;
        10'b0000000100 : logsin1 = mux_in_sin4;
        10'b0000000101 : logsin1 = mux_in_sin5;
        10'b0000000110 : logsin1 = mux_in_sin6;
        10'b0000000111 : logsin1 = mux_in_sin7;
        10'b0000001000 : logsin1 = mux_in_sin8;
        10'b0000001001 : logsin1 = mux_in_sin9;
        10'b0000001010 : logsin1 = mux_in_sin10;
        10'b0000001011 : logsin1 = mux_in_sin11;
        10'b0000001100 : logsin1 = mux_in_sin12;
        10'b0000001101 : logsin1 = mux_in_sin13;
        10'b0000001110 : logsin1 = mux_in_sin14;
        10'b0000001111 : logsin1 = mux_in_sin15;
        10'b0000010000 : logsin1 = mux_in_sin16;
        10'b0000010001 : logsin1 = mux_in_sin17;
        10'b0000010010 : logsin1 = mux_in_sin18;
        10'b0000010011 : logsin1 = mux_in_sin19;
        10'b0000010100 : logsin1 = mux_in_sin20;
        10'b0000010101 : logsin1 = mux_in_sin21;
        10'b0000010110 : logsin1 = mux_in_sin22;
        10'b0000010111 : logsin1 = mux_in_sin23;
        10'b0000011000 : logsin1 = mux_in_sin24;
        10'b0000011001 : logsin1 = mux_in_sin25;
        10'b0000011010 : logsin1 = mux_in_sin26;
        10'b0000011011 : logsin1 = mux_in_sin27;
        10'b0000011100 : logsin1 = mux_in_sin28;
        10'b0000011101 : logsin1 = mux_in_sin29;
        10'b0000011110 : logsin1 = mux_in_sin30;
        10'b0000011111 : logsin1 = mux_in_sin31;
        10'b0000100000 : logsin1 = mux_in_sin32;
        10'b0000100001 : logsin1 = mux_in_sin33;
        10'b0000100010 : logsin1 = mux_in_sin34;
        10'b0000100011 : logsin1 = mux_in_sin35;
        10'b0000100100 : logsin1 = mux_in_sin36;
        10'b0000100101 : logsin1 = mux_in_sin37;
        10'b0000100110 : logsin1 = mux_in_sin38;
        10'b0000100111 : logsin1 = mux_in_sin39;
        10'b0000101000 : logsin1 = mux_in_sin40;
        10'b0000101001 : logsin1 = mux_in_sin41;
        10'b0000101010 : logsin1 = mux_in_sin42;
        10'b0000101011 : logsin1 = mux_in_sin43;
        10'b0000101100 : logsin1 = mux_in_sin44;
        10'b0000101101 : logsin1 = mux_in_sin45;
        10'b0000101110 : logsin1 = mux_in_sin46;
        10'b0000101111 : logsin1 = mux_in_sin47;
        10'b0000110000 : logsin1 = mux_in_sin48;
        10'b0000110001 : logsin1 = mux_in_sin49;
        10'b0000110010 : logsin1 = mux_in_sin50;
        10'b0000110011 : logsin1 = mux_in_sin51;
        10'b0000110100 : logsin1 = mux_in_sin52;
        10'b0000110101 : logsin1 = mux_in_sin53;
        10'b0000110110 : logsin1 = mux_in_sin54;
        10'b0000110111 : logsin1 = mux_in_sin55;
        10'b0000111000 : logsin1 = mux_in_sin56;
        10'b0000111001 : logsin1 = mux_in_sin57;
        10'b0000111010 : logsin1 = mux_in_sin58;
        10'b0000111011 : logsin1 = mux_in_sin59;
        10'b0000111100 : logsin1 = mux_in_sin60;
        10'b0000111101 : logsin1 = mux_in_sin61;
        10'b0000111110 : logsin1 = mux_in_sin62;
        10'b0000111111 : logsin1 = mux_in_sin63;
        10'b0001000000 : logsin1 = mux_in_sin64;
        10'b0001000001 : logsin1 = mux_in_sin65;
        10'b0001000010 : logsin1 = mux_in_sin66;
        10'b0001000011 : logsin1 = mux_in_sin67;
        10'b0001000100 : logsin1 = mux_in_sin68;
        10'b0001000101 : logsin1 = mux_in_sin69;
        10'b0001000110 : logsin1 = mux_in_sin70;
        10'b0001000111 : logsin1 = mux_in_sin71;
        10'b0001001000 : logsin1 = mux_in_sin72;
        10'b0001001001 : logsin1 = mux_in_sin73;
        10'b0001001010 : logsin1 = mux_in_sin74;
        10'b0001001011 : logsin1 = mux_in_sin75;
        10'b0001001100 : logsin1 = mux_in_sin76;
        10'b0001001101 : logsin1 = mux_in_sin77;
        10'b0001001110 : logsin1 = mux_in_sin78;
        10'b0001001111 : logsin1 = mux_in_sin79;
        10'b0001010000 : logsin1 = mux_in_sin80;
        10'b0001010001 : logsin1 = mux_in_sin81;
        10'b0001010010 : logsin1 = mux_in_sin82;
        10'b0001010011 : logsin1 = mux_in_sin83;
        10'b0001010100 : logsin1 = mux_in_sin84;
        10'b0001010101 : logsin1 = mux_in_sin85;
        10'b0001010110 : logsin1 = mux_in_sin86;
        10'b0001010111 : logsin1 = mux_in_sin87;
        10'b0001011000 : logsin1 = mux_in_sin88;
        10'b0001011001 : logsin1 = mux_in_sin89;
        10'b0001011010 : logsin1 = mux_in_sin90;
        10'b0001011011 : logsin1 = mux_in_sin91;
        10'b0001011100 : logsin1 = mux_in_sin92;
        10'b0001011101 : logsin1 = mux_in_sin93;
        10'b0001011110 : logsin1 = mux_in_sin94;
        10'b0001011111 : logsin1 = mux_in_sin95;
        10'b0001100000 : logsin1 = mux_in_sin96;
        10'b0001100001 : logsin1 = mux_in_sin97;
        10'b0001100010 : logsin1 = mux_in_sin98;
        10'b0001100011 : logsin1 = mux_in_sin99;
        10'b0001100100 : logsin1 = mux_in_sin100;
        10'b0001100101 : logsin1 = mux_in_sin101;
        10'b0001100110 : logsin1 = mux_in_sin102;
        10'b0001100111 : logsin1 = mux_in_sin103;
        10'b0001101000 : logsin1 = mux_in_sin104;
        10'b0001101001 : logsin1 = mux_in_sin105;
        10'b0001101010 : logsin1 = mux_in_sin106;
        10'b0001101011 : logsin1 = mux_in_sin107;
        10'b0001101100 : logsin1 = mux_in_sin108;
        10'b0001101101 : logsin1 = mux_in_sin109;
        10'b0001101110 : logsin1 = mux_in_sin110;
        10'b0001101111 : logsin1 = mux_in_sin111;
        10'b0001110000 : logsin1 = mux_in_sin112;
        10'b0001110001 : logsin1 = mux_in_sin113;
        10'b0001110010 : logsin1 = mux_in_sin114;
        10'b0001110011 : logsin1 = mux_in_sin115;
        10'b0001110100 : logsin1 = mux_in_sin116;
        10'b0001110101 : logsin1 = mux_in_sin117;
        10'b0001110110 : logsin1 = mux_in_sin118;
        10'b0001110111 : logsin1 = mux_in_sin119;
        10'b0001111000 : logsin1 = mux_in_sin120;
        10'b0001111001 : logsin1 = mux_in_sin121;
        10'b0001111010 : logsin1 = mux_in_sin122;
        10'b0001111011 : logsin1 = mux_in_sin123;
        10'b0001111100 : logsin1 = mux_in_sin124;
        10'b0001111101 : logsin1 = mux_in_sin125;
        10'b0001111110 : logsin1 = mux_in_sin126;
        10'b0001111111 : logsin1 = mux_in_sin127;
        10'b0010000000 : logsin1 = mux_in_sin128;
        10'b0010000001 : logsin1 = mux_in_sin129;
        10'b0010000010 : logsin1 = mux_in_sin130;
        10'b0010000011 : logsin1 = mux_in_sin131;
        10'b0010000100 : logsin1 = mux_in_sin132;
        10'b0010000101 : logsin1 = mux_in_sin133;
        10'b0010000110 : logsin1 = mux_in_sin134;
        10'b0010000111 : logsin1 = mux_in_sin135;
        10'b0010001000 : logsin1 = mux_in_sin136;
        10'b0010001001 : logsin1 = mux_in_sin137;
        10'b0010001010 : logsin1 = mux_in_sin138;
        10'b0010001011 : logsin1 = mux_in_sin139;
        10'b0010001100 : logsin1 = mux_in_sin140;
        10'b0010001101 : logsin1 = mux_in_sin141;
        10'b0010001110 : logsin1 = mux_in_sin142;
        10'b0010001111 : logsin1 = mux_in_sin143;
        10'b0010010000 : logsin1 = mux_in_sin144;
        10'b0010010001 : logsin1 = mux_in_sin145;
        10'b0010010010 : logsin1 = mux_in_sin146;
        10'b0010010011 : logsin1 = mux_in_sin147;
        10'b0010010100 : logsin1 = mux_in_sin148;
        10'b0010010101 : logsin1 = mux_in_sin149;
        10'b0010010110 : logsin1 = mux_in_sin150;
        10'b0010010111 : logsin1 = mux_in_sin151;
        10'b0010011000 : logsin1 = mux_in_sin152;
        10'b0010011001 : logsin1 = mux_in_sin153;
        10'b0010011010 : logsin1 = mux_in_sin154;
        10'b0010011011 : logsin1 = mux_in_sin155;
        10'b0010011100 : logsin1 = mux_in_sin156;
        10'b0010011101 : logsin1 = mux_in_sin157;
        10'b0010011110 : logsin1 = mux_in_sin158;
        10'b0010011111 : logsin1 = mux_in_sin159;
        10'b0010100000 : logsin1 = mux_in_sin160;
        10'b0010100001 : logsin1 = mux_in_sin161;
        10'b0010100010 : logsin1 = mux_in_sin162;
        10'b0010100011 : logsin1 = mux_in_sin163;
        10'b0010100100 : logsin1 = mux_in_sin164;
        10'b0010100101 : logsin1 = mux_in_sin165;
        10'b0010100110 : logsin1 = mux_in_sin166;
        10'b0010100111 : logsin1 = mux_in_sin167;
        10'b0010101000 : logsin1 = mux_in_sin168;
        10'b0010101001 : logsin1 = mux_in_sin169;
        10'b0010101010 : logsin1 = mux_in_sin170;
        10'b0010101011 : logsin1 = mux_in_sin171;
        10'b0010101100 : logsin1 = mux_in_sin172;
        10'b0010101101 : logsin1 = mux_in_sin173;
        10'b0010101110 : logsin1 = mux_in_sin174;
        10'b0010101111 : logsin1 = mux_in_sin175;
        10'b0010110000 : logsin1 = mux_in_sin176;
        10'b0010110001 : logsin1 = mux_in_sin177;
        10'b0010110010 : logsin1 = mux_in_sin178;
        10'b0010110011 : logsin1 = mux_in_sin179;
        10'b0010110100 : logsin1 = mux_in_sin180;
        10'b0010110101 : logsin1 = mux_in_sin181;
        10'b0010110110 : logsin1 = mux_in_sin182;
        10'b0010110111 : logsin1 = mux_in_sin183;
        10'b0010111000 : logsin1 = mux_in_sin184;
        10'b0010111001 : logsin1 = mux_in_sin185;
        10'b0010111010 : logsin1 = mux_in_sin186;
        10'b0010111011 : logsin1 = mux_in_sin187;
        10'b0010111100 : logsin1 = mux_in_sin188;
        10'b0010111101 : logsin1 = mux_in_sin189;
        10'b0010111110 : logsin1 = mux_in_sin190;
        10'b0010111111 : logsin1 = mux_in_sin191;
        10'b0011000000 : logsin1 = mux_in_sin192;
        10'b0011000001 : logsin1 = mux_in_sin193;
        10'b0011000010 : logsin1 = mux_in_sin194;
        10'b0011000011 : logsin1 = mux_in_sin195;
        10'b0011000100 : logsin1 = mux_in_sin196;
        10'b0011000101 : logsin1 = mux_in_sin197;
        10'b0011000110 : logsin1 = mux_in_sin198;
        10'b0011000111 : logsin1 = mux_in_sin199;
        10'b0011001000 : logsin1 = mux_in_sin200;
        10'b0011001001 : logsin1 = mux_in_sin201;
        10'b0011001010 : logsin1 = mux_in_sin202;
        10'b0011001011 : logsin1 = mux_in_sin203;
        10'b0011001100 : logsin1 = mux_in_sin204;
        10'b0011001101 : logsin1 = mux_in_sin205;
        10'b0011001110 : logsin1 = mux_in_sin206;
        10'b0011001111 : logsin1 = mux_in_sin207;
        10'b0011010000 : logsin1 = mux_in_sin208;
        10'b0011010001 : logsin1 = mux_in_sin209;
        10'b0011010010 : logsin1 = mux_in_sin210;
        10'b0011010011 : logsin1 = mux_in_sin211;
        10'b0011010100 : logsin1 = mux_in_sin212;
        10'b0011010101 : logsin1 = mux_in_sin213;
        10'b0011010110 : logsin1 = mux_in_sin214;
        10'b0011010111 : logsin1 = mux_in_sin215;
        10'b0011011000 : logsin1 = mux_in_sin216;
        10'b0011011001 : logsin1 = mux_in_sin217;
        10'b0011011010 : logsin1 = mux_in_sin218;
        10'b0011011011 : logsin1 = mux_in_sin219;
        10'b0011011100 : logsin1 = mux_in_sin220;
        10'b0011011101 : logsin1 = mux_in_sin221;
        10'b0011011110 : logsin1 = mux_in_sin222;
        10'b0011011111 : logsin1 = mux_in_sin223;
        10'b0011100000 : logsin1 = mux_in_sin224;
        10'b0011100001 : logsin1 = mux_in_sin225;
        10'b0011100010 : logsin1 = mux_in_sin226;
        10'b0011100011 : logsin1 = mux_in_sin227;
        10'b0011100100 : logsin1 = mux_in_sin228;
        10'b0011100101 : logsin1 = mux_in_sin229;
        10'b0011100110 : logsin1 = mux_in_sin230;
        10'b0011100111 : logsin1 = mux_in_sin231;
        10'b0011101000 : logsin1 = mux_in_sin232;
        10'b0011101001 : logsin1 = mux_in_sin233;
        10'b0011101010 : logsin1 = mux_in_sin234;
        10'b0011101011 : logsin1 = mux_in_sin235;
        10'b0011101100 : logsin1 = mux_in_sin236;
        10'b0011101101 : logsin1 = mux_in_sin237;
        10'b0011101110 : logsin1 = mux_in_sin238;
        10'b0011101111 : logsin1 = mux_in_sin239;
        10'b0011110000 : logsin1 = mux_in_sin240;
        10'b0011110001 : logsin1 = mux_in_sin241;
        10'b0011110010 : logsin1 = mux_in_sin242;
        10'b0011110011 : logsin1 = mux_in_sin243;
        10'b0011110100 : logsin1 = mux_in_sin244;
        10'b0011110101 : logsin1 = mux_in_sin245;
        10'b0011110110 : logsin1 = mux_in_sin246;
        10'b0011110111 : logsin1 = mux_in_sin247;
        10'b0011111000 : logsin1 = mux_in_sin248;
        10'b0011111001 : logsin1 = mux_in_sin249;
        10'b0011111010 : logsin1 = mux_in_sin250;
        10'b0011111011 : logsin1 = mux_in_sin251;
        10'b0011111100 : logsin1 = mux_in_sin252;
        10'b0011111101 : logsin1 = mux_in_sin253;
        10'b0011111110 : logsin1 = mux_in_sin254;
        10'b0011111111 : logsin1 = mux_in_sin255;
        10'b0100000000 : logsin1 = mux_in_sin256;
        10'b0100000001 : logsin1 = mux_in_sin257;
        10'b0100000010 : logsin1 = mux_in_sin258;
        10'b0100000011 : logsin1 = mux_in_sin259;
        10'b0100000100 : logsin1 = mux_in_sin260;
        10'b0100000101 : logsin1 = mux_in_sin261;
        10'b0100000110 : logsin1 = mux_in_sin262;
        10'b0100000111 : logsin1 = mux_in_sin263;
        10'b0100001000 : logsin1 = mux_in_sin264;
        10'b0100001001 : logsin1 = mux_in_sin265;
        10'b0100001010 : logsin1 = mux_in_sin266;
        10'b0100001011 : logsin1 = mux_in_sin267;
        10'b0100001100 : logsin1 = mux_in_sin268;
        10'b0100001101 : logsin1 = mux_in_sin269;
        10'b0100001110 : logsin1 = mux_in_sin270;
        10'b0100001111 : logsin1 = mux_in_sin271;
        10'b0100010000 : logsin1 = mux_in_sin272;
        10'b0100010001 : logsin1 = mux_in_sin273;
        10'b0100010010 : logsin1 = mux_in_sin274;
        10'b0100010011 : logsin1 = mux_in_sin275;
        10'b0100010100 : logsin1 = mux_in_sin276;
        10'b0100010101 : logsin1 = mux_in_sin277;
        10'b0100010110 : logsin1 = mux_in_sin278;
        10'b0100010111 : logsin1 = mux_in_sin279;
        10'b0100011000 : logsin1 = mux_in_sin280;
        10'b0100011001 : logsin1 = mux_in_sin281;
        10'b0100011010 : logsin1 = mux_in_sin282;
        10'b0100011011 : logsin1 = mux_in_sin283;
        10'b0100011100 : logsin1 = mux_in_sin284;
        10'b0100011101 : logsin1 = mux_in_sin285;
        10'b0100011110 : logsin1 = mux_in_sin286;
        10'b0100011111 : logsin1 = mux_in_sin287;
        10'b0100100000 : logsin1 = mux_in_sin288;
        10'b0100100001 : logsin1 = mux_in_sin289;
        10'b0100100010 : logsin1 = mux_in_sin290;
        10'b0100100011 : logsin1 = mux_in_sin291;
        10'b0100100100 : logsin1 = mux_in_sin292;
        10'b0100100101 : logsin1 = mux_in_sin293;
        10'b0100100110 : logsin1 = mux_in_sin294;
        10'b0100100111 : logsin1 = mux_in_sin295;
        10'b0100101000 : logsin1 = mux_in_sin296;
        10'b0100101001 : logsin1 = mux_in_sin297;
        10'b0100101010 : logsin1 = mux_in_sin298;
        10'b0100101011 : logsin1 = mux_in_sin299;
        10'b0100101100 : logsin1 = mux_in_sin300;
        10'b0100101101 : logsin1 = mux_in_sin301;
        10'b0100101110 : logsin1 = mux_in_sin302;
        10'b0100101111 : logsin1 = mux_in_sin303;
        10'b0100110000 : logsin1 = mux_in_sin304;
        10'b0100110001 : logsin1 = mux_in_sin305;
        10'b0100110010 : logsin1 = mux_in_sin306;
        10'b0100110011 : logsin1 = mux_in_sin307;
        10'b0100110100 : logsin1 = mux_in_sin308;
        10'b0100110101 : logsin1 = mux_in_sin309;
        10'b0100110110 : logsin1 = mux_in_sin310;
        10'b0100110111 : logsin1 = mux_in_sin311;
        10'b0100111000 : logsin1 = mux_in_sin312;
        10'b0100111001 : logsin1 = mux_in_sin313;
        10'b0100111010 : logsin1 = mux_in_sin314;
        10'b0100111011 : logsin1 = mux_in_sin315;
        10'b0100111100 : logsin1 = mux_in_sin316;
        10'b0100111101 : logsin1 = mux_in_sin317;
        10'b0100111110 : logsin1 = mux_in_sin318;
        10'b0100111111 : logsin1 = mux_in_sin319;
        10'b0101000000 : logsin1 = mux_in_sin320;
        10'b0101000001 : logsin1 = mux_in_sin321;
        10'b0101000010 : logsin1 = mux_in_sin322;
        10'b0101000011 : logsin1 = mux_in_sin323;
        10'b0101000100 : logsin1 = mux_in_sin324;
        10'b0101000101 : logsin1 = mux_in_sin325;
        10'b0101000110 : logsin1 = mux_in_sin326;
        10'b0101000111 : logsin1 = mux_in_sin327;
        10'b0101001000 : logsin1 = mux_in_sin328;
        10'b0101001001 : logsin1 = mux_in_sin329;
        10'b0101001010 : logsin1 = mux_in_sin330;
        10'b0101001011 : logsin1 = mux_in_sin331;
        10'b0101001100 : logsin1 = mux_in_sin332;
        10'b0101001101 : logsin1 = mux_in_sin333;
        10'b0101001110 : logsin1 = mux_in_sin334;
        10'b0101001111 : logsin1 = mux_in_sin335;
        10'b0101010000 : logsin1 = mux_in_sin336;
        10'b0101010001 : logsin1 = mux_in_sin337;
        10'b0101010010 : logsin1 = mux_in_sin338;
        10'b0101010011 : logsin1 = mux_in_sin339;
        10'b0101010100 : logsin1 = mux_in_sin340;
        10'b0101010101 : logsin1 = mux_in_sin341;
        10'b0101010110 : logsin1 = mux_in_sin342;
        10'b0101010111 : logsin1 = mux_in_sin343;
        10'b0101011000 : logsin1 = mux_in_sin344;
        10'b0101011001 : logsin1 = mux_in_sin345;
        10'b0101011010 : logsin1 = mux_in_sin346;
        10'b0101011011 : logsin1 = mux_in_sin347;
        10'b0101011100 : logsin1 = mux_in_sin348;
        10'b0101011101 : logsin1 = mux_in_sin349;
        10'b0101011110 : logsin1 = mux_in_sin350;
        10'b0101011111 : logsin1 = mux_in_sin351;
        10'b0101100000 : logsin1 = mux_in_sin352;
        10'b0101100001 : logsin1 = mux_in_sin353;
        10'b0101100010 : logsin1 = mux_in_sin354;
        10'b0101100011 : logsin1 = mux_in_sin355;
        10'b0101100100 : logsin1 = mux_in_sin356;
        10'b0101100101 : logsin1 = mux_in_sin357;
        10'b0101100110 : logsin1 = mux_in_sin358;
        10'b0101100111 : logsin1 = mux_in_sin359;
        10'b0101101000 : logsin1 = mux_in_sin360;
        10'b0101101001 : logsin1 = mux_in_sin361;
        10'b0101101010 : logsin1 = mux_in_sin362;
        10'b0101101011 : logsin1 = mux_in_sin363;
        10'b0101101100 : logsin1 = mux_in_sin364;
        10'b0101101101 : logsin1 = mux_in_sin365;
        10'b0101101110 : logsin1 = mux_in_sin366;
        10'b0101101111 : logsin1 = mux_in_sin367;
        10'b0101110000 : logsin1 = mux_in_sin368;
        10'b0101110001 : logsin1 = mux_in_sin369;
        10'b0101110010 : logsin1 = mux_in_sin370;
        10'b0101110011 : logsin1 = mux_in_sin371;
        10'b0101110100 : logsin1 = mux_in_sin372;
        10'b0101110101 : logsin1 = mux_in_sin373;
        10'b0101110110 : logsin1 = mux_in_sin374;
        10'b0101110111 : logsin1 = mux_in_sin375;
        10'b0101111000 : logsin1 = mux_in_sin376;
        10'b0101111001 : logsin1 = mux_in_sin377;
        10'b0101111010 : logsin1 = mux_in_sin378;
        10'b0101111011 : logsin1 = mux_in_sin379;
        10'b0101111100 : logsin1 = mux_in_sin380;
        10'b0101111101 : logsin1 = mux_in_sin381;
        10'b0101111110 : logsin1 = mux_in_sin382;
        10'b0101111111 : logsin1 = mux_in_sin383;
        10'b0110000000 : logsin1 = mux_in_sin384;
        10'b0110000001 : logsin1 = mux_in_sin385;
        10'b0110000010 : logsin1 = mux_in_sin386;
        10'b0110000011 : logsin1 = mux_in_sin387;
        10'b0110000100 : logsin1 = mux_in_sin388;
        10'b0110000101 : logsin1 = mux_in_sin389;
        10'b0110000110 : logsin1 = mux_in_sin390;
        10'b0110000111 : logsin1 = mux_in_sin391;
        10'b0110001000 : logsin1 = mux_in_sin392;
        10'b0110001001 : logsin1 = mux_in_sin393;
        10'b0110001010 : logsin1 = mux_in_sin394;
        10'b0110001011 : logsin1 = mux_in_sin395;
        10'b0110001100 : logsin1 = mux_in_sin396;
        10'b0110001101 : logsin1 = mux_in_sin397;
        10'b0110001110 : logsin1 = mux_in_sin398;
        10'b0110001111 : logsin1 = mux_in_sin399;
        10'b0110010000 : logsin1 = mux_in_sin400;
        10'b0110010001 : logsin1 = mux_in_sin401;
        10'b0110010010 : logsin1 = mux_in_sin402;
        10'b0110010011 : logsin1 = mux_in_sin403;
        10'b0110010100 : logsin1 = mux_in_sin404;
        10'b0110010101 : logsin1 = mux_in_sin405;
        10'b0110010110 : logsin1 = mux_in_sin406;
        10'b0110010111 : logsin1 = mux_in_sin407;
        10'b0110011000 : logsin1 = mux_in_sin408;
        10'b0110011001 : logsin1 = mux_in_sin409;
        10'b0110011010 : logsin1 = mux_in_sin410;
        10'b0110011011 : logsin1 = mux_in_sin411;
        10'b0110011100 : logsin1 = mux_in_sin412;
        10'b0110011101 : logsin1 = mux_in_sin413;
        10'b0110011110 : logsin1 = mux_in_sin414;
        10'b0110011111 : logsin1 = mux_in_sin415;
        10'b0110100000 : logsin1 = mux_in_sin416;
        10'b0110100001 : logsin1 = mux_in_sin417;
        10'b0110100010 : logsin1 = mux_in_sin418;
        10'b0110100011 : logsin1 = mux_in_sin419;
        10'b0110100100 : logsin1 = mux_in_sin420;
        10'b0110100101 : logsin1 = mux_in_sin421;
        10'b0110100110 : logsin1 = mux_in_sin422;
        10'b0110100111 : logsin1 = mux_in_sin423;
        10'b0110101000 : logsin1 = mux_in_sin424;
        10'b0110101001 : logsin1 = mux_in_sin425;
        10'b0110101010 : logsin1 = mux_in_sin426;
        10'b0110101011 : logsin1 = mux_in_sin427;
        10'b0110101100 : logsin1 = mux_in_sin428;
        10'b0110101101 : logsin1 = mux_in_sin429;
        10'b0110101110 : logsin1 = mux_in_sin430;
        10'b0110101111 : logsin1 = mux_in_sin431;
        10'b0110110000 : logsin1 = mux_in_sin432;
        10'b0110110001 : logsin1 = mux_in_sin433;
        10'b0110110010 : logsin1 = mux_in_sin434;
        10'b0110110011 : logsin1 = mux_in_sin435;
        10'b0110110100 : logsin1 = mux_in_sin436;
        10'b0110110101 : logsin1 = mux_in_sin437;
        10'b0110110110 : logsin1 = mux_in_sin438;
        10'b0110110111 : logsin1 = mux_in_sin439;
        10'b0110111000 : logsin1 = mux_in_sin440;
        10'b0110111001 : logsin1 = mux_in_sin441;
        10'b0110111010 : logsin1 = mux_in_sin442;
        10'b0110111011 : logsin1 = mux_in_sin443;
        10'b0110111100 : logsin1 = mux_in_sin444;
        10'b0110111101 : logsin1 = mux_in_sin445;
        10'b0110111110 : logsin1 = mux_in_sin446;
        10'b0110111111 : logsin1 = mux_in_sin447;
        10'b0111000000 : logsin1 = mux_in_sin448;
        10'b0111000001 : logsin1 = mux_in_sin449;
        10'b0111000010 : logsin1 = mux_in_sin450;
        10'b0111000011 : logsin1 = mux_in_sin451;
        10'b0111000100 : logsin1 = mux_in_sin452;
        10'b0111000101 : logsin1 = mux_in_sin453;
        10'b0111000110 : logsin1 = mux_in_sin454;
        10'b0111000111 : logsin1 = mux_in_sin455;
        10'b0111001000 : logsin1 = mux_in_sin456;
        10'b0111001001 : logsin1 = mux_in_sin457;
        10'b0111001010 : logsin1 = mux_in_sin458;
        10'b0111001011 : logsin1 = mux_in_sin459;
        10'b0111001100 : logsin1 = mux_in_sin460;
        10'b0111001101 : logsin1 = mux_in_sin461;
        10'b0111001110 : logsin1 = mux_in_sin462;
        10'b0111001111 : logsin1 = mux_in_sin463;
        10'b0111010000 : logsin1 = mux_in_sin464;
        10'b0111010001 : logsin1 = mux_in_sin465;
        10'b0111010010 : logsin1 = mux_in_sin466;
        10'b0111010011 : logsin1 = mux_in_sin467;
        10'b0111010100 : logsin1 = mux_in_sin468;
        10'b0111010101 : logsin1 = mux_in_sin469;
        10'b0111010110 : logsin1 = mux_in_sin470;
        10'b0111010111 : logsin1 = mux_in_sin471;
        10'b0111011000 : logsin1 = mux_in_sin472;
        10'b0111011001 : logsin1 = mux_in_sin473;
        10'b0111011010 : logsin1 = mux_in_sin474;
        10'b0111011011 : logsin1 = mux_in_sin475;
        10'b0111011100 : logsin1 = mux_in_sin476;
        10'b0111011101 : logsin1 = mux_in_sin477;
        10'b0111011110 : logsin1 = mux_in_sin478;
        10'b0111011111 : logsin1 = mux_in_sin479;
        10'b0111100000 : logsin1 = mux_in_sin480;
        10'b0111100001 : logsin1 = mux_in_sin481;
        10'b0111100010 : logsin1 = mux_in_sin482;
        10'b0111100011 : logsin1 = mux_in_sin483;
        10'b0111100100 : logsin1 = mux_in_sin484;
        10'b0111100101 : logsin1 = mux_in_sin485;
        10'b0111100110 : logsin1 = mux_in_sin486;
        10'b0111100111 : logsin1 = mux_in_sin487;
        10'b0111101000 : logsin1 = mux_in_sin488;
        10'b0111101001 : logsin1 = mux_in_sin489;
        10'b0111101010 : logsin1 = mux_in_sin490;
        10'b0111101011 : logsin1 = mux_in_sin491;
        10'b0111101100 : logsin1 = mux_in_sin492;
        10'b0111101101 : logsin1 = mux_in_sin493;
        10'b0111101110 : logsin1 = mux_in_sin494;
        10'b0111101111 : logsin1 = mux_in_sin495;
        10'b0111110000 : logsin1 = mux_in_sin496;
        10'b0111110001 : logsin1 = mux_in_sin497;
        10'b0111110010 : logsin1 = mux_in_sin498;
        10'b0111110011 : logsin1 = mux_in_sin499;
        10'b0111110100 : logsin1 = mux_in_sin500;
        10'b0111110101 : logsin1 = mux_in_sin501;
        10'b0111110110 : logsin1 = mux_in_sin502;
        10'b0111110111 : logsin1 = mux_in_sin503;
        10'b0111111000 : logsin1 = mux_in_sin504;
        10'b0111111001 : logsin1 = mux_in_sin505;
        10'b0111111010 : logsin1 = mux_in_sin506;
        10'b0111111011 : logsin1 = mux_in_sin507;
        10'b0111111100 : logsin1 = mux_in_sin508;
        10'b0111111101 : logsin1 = mux_in_sin509;
        10'b0111111110 : logsin1 = mux_in_sin510;
        10'b0111111111 : logsin1 = mux_in_sin511;
        10'b1000000000 : logsin1 = mux_in_sin512;
        default: logsin1 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in2)
        10'b0000000000 : logsin2 = mux_in_sin0;
        10'b0000000001 : logsin2 = mux_in_sin1;
        10'b0000000010 : logsin2 = mux_in_sin2;
        10'b0000000011 : logsin2 = mux_in_sin3;
        10'b0000000100 : logsin2 = mux_in_sin4;
        10'b0000000101 : logsin2 = mux_in_sin5;
        10'b0000000110 : logsin2 = mux_in_sin6;
        10'b0000000111 : logsin2 = mux_in_sin7;
        10'b0000001000 : logsin2 = mux_in_sin8;
        10'b0000001001 : logsin2 = mux_in_sin9;
        10'b0000001010 : logsin2 = mux_in_sin10;
        10'b0000001011 : logsin2 = mux_in_sin11;
        10'b0000001100 : logsin2 = mux_in_sin12;
        10'b0000001101 : logsin2 = mux_in_sin13;
        10'b0000001110 : logsin2 = mux_in_sin14;
        10'b0000001111 : logsin2 = mux_in_sin15;
        10'b0000010000 : logsin2 = mux_in_sin16;
        10'b0000010001 : logsin2 = mux_in_sin17;
        10'b0000010010 : logsin2 = mux_in_sin18;
        10'b0000010011 : logsin2 = mux_in_sin19;
        10'b0000010100 : logsin2 = mux_in_sin20;
        10'b0000010101 : logsin2 = mux_in_sin21;
        10'b0000010110 : logsin2 = mux_in_sin22;
        10'b0000010111 : logsin2 = mux_in_sin23;
        10'b0000011000 : logsin2 = mux_in_sin24;
        10'b0000011001 : logsin2 = mux_in_sin25;
        10'b0000011010 : logsin2 = mux_in_sin26;
        10'b0000011011 : logsin2 = mux_in_sin27;
        10'b0000011100 : logsin2 = mux_in_sin28;
        10'b0000011101 : logsin2 = mux_in_sin29;
        10'b0000011110 : logsin2 = mux_in_sin30;
        10'b0000011111 : logsin2 = mux_in_sin31;
        10'b0000100000 : logsin2 = mux_in_sin32;
        10'b0000100001 : logsin2 = mux_in_sin33;
        10'b0000100010 : logsin2 = mux_in_sin34;
        10'b0000100011 : logsin2 = mux_in_sin35;
        10'b0000100100 : logsin2 = mux_in_sin36;
        10'b0000100101 : logsin2 = mux_in_sin37;
        10'b0000100110 : logsin2 = mux_in_sin38;
        10'b0000100111 : logsin2 = mux_in_sin39;
        10'b0000101000 : logsin2 = mux_in_sin40;
        10'b0000101001 : logsin2 = mux_in_sin41;
        10'b0000101010 : logsin2 = mux_in_sin42;
        10'b0000101011 : logsin2 = mux_in_sin43;
        10'b0000101100 : logsin2 = mux_in_sin44;
        10'b0000101101 : logsin2 = mux_in_sin45;
        10'b0000101110 : logsin2 = mux_in_sin46;
        10'b0000101111 : logsin2 = mux_in_sin47;
        10'b0000110000 : logsin2 = mux_in_sin48;
        10'b0000110001 : logsin2 = mux_in_sin49;
        10'b0000110010 : logsin2 = mux_in_sin50;
        10'b0000110011 : logsin2 = mux_in_sin51;
        10'b0000110100 : logsin2 = mux_in_sin52;
        10'b0000110101 : logsin2 = mux_in_sin53;
        10'b0000110110 : logsin2 = mux_in_sin54;
        10'b0000110111 : logsin2 = mux_in_sin55;
        10'b0000111000 : logsin2 = mux_in_sin56;
        10'b0000111001 : logsin2 = mux_in_sin57;
        10'b0000111010 : logsin2 = mux_in_sin58;
        10'b0000111011 : logsin2 = mux_in_sin59;
        10'b0000111100 : logsin2 = mux_in_sin60;
        10'b0000111101 : logsin2 = mux_in_sin61;
        10'b0000111110 : logsin2 = mux_in_sin62;
        10'b0000111111 : logsin2 = mux_in_sin63;
        10'b0001000000 : logsin2 = mux_in_sin64;
        10'b0001000001 : logsin2 = mux_in_sin65;
        10'b0001000010 : logsin2 = mux_in_sin66;
        10'b0001000011 : logsin2 = mux_in_sin67;
        10'b0001000100 : logsin2 = mux_in_sin68;
        10'b0001000101 : logsin2 = mux_in_sin69;
        10'b0001000110 : logsin2 = mux_in_sin70;
        10'b0001000111 : logsin2 = mux_in_sin71;
        10'b0001001000 : logsin2 = mux_in_sin72;
        10'b0001001001 : logsin2 = mux_in_sin73;
        10'b0001001010 : logsin2 = mux_in_sin74;
        10'b0001001011 : logsin2 = mux_in_sin75;
        10'b0001001100 : logsin2 = mux_in_sin76;
        10'b0001001101 : logsin2 = mux_in_sin77;
        10'b0001001110 : logsin2 = mux_in_sin78;
        10'b0001001111 : logsin2 = mux_in_sin79;
        10'b0001010000 : logsin2 = mux_in_sin80;
        10'b0001010001 : logsin2 = mux_in_sin81;
        10'b0001010010 : logsin2 = mux_in_sin82;
        10'b0001010011 : logsin2 = mux_in_sin83;
        10'b0001010100 : logsin2 = mux_in_sin84;
        10'b0001010101 : logsin2 = mux_in_sin85;
        10'b0001010110 : logsin2 = mux_in_sin86;
        10'b0001010111 : logsin2 = mux_in_sin87;
        10'b0001011000 : logsin2 = mux_in_sin88;
        10'b0001011001 : logsin2 = mux_in_sin89;
        10'b0001011010 : logsin2 = mux_in_sin90;
        10'b0001011011 : logsin2 = mux_in_sin91;
        10'b0001011100 : logsin2 = mux_in_sin92;
        10'b0001011101 : logsin2 = mux_in_sin93;
        10'b0001011110 : logsin2 = mux_in_sin94;
        10'b0001011111 : logsin2 = mux_in_sin95;
        10'b0001100000 : logsin2 = mux_in_sin96;
        10'b0001100001 : logsin2 = mux_in_sin97;
        10'b0001100010 : logsin2 = mux_in_sin98;
        10'b0001100011 : logsin2 = mux_in_sin99;
        10'b0001100100 : logsin2 = mux_in_sin100;
        10'b0001100101 : logsin2 = mux_in_sin101;
        10'b0001100110 : logsin2 = mux_in_sin102;
        10'b0001100111 : logsin2 = mux_in_sin103;
        10'b0001101000 : logsin2 = mux_in_sin104;
        10'b0001101001 : logsin2 = mux_in_sin105;
        10'b0001101010 : logsin2 = mux_in_sin106;
        10'b0001101011 : logsin2 = mux_in_sin107;
        10'b0001101100 : logsin2 = mux_in_sin108;
        10'b0001101101 : logsin2 = mux_in_sin109;
        10'b0001101110 : logsin2 = mux_in_sin110;
        10'b0001101111 : logsin2 = mux_in_sin111;
        10'b0001110000 : logsin2 = mux_in_sin112;
        10'b0001110001 : logsin2 = mux_in_sin113;
        10'b0001110010 : logsin2 = mux_in_sin114;
        10'b0001110011 : logsin2 = mux_in_sin115;
        10'b0001110100 : logsin2 = mux_in_sin116;
        10'b0001110101 : logsin2 = mux_in_sin117;
        10'b0001110110 : logsin2 = mux_in_sin118;
        10'b0001110111 : logsin2 = mux_in_sin119;
        10'b0001111000 : logsin2 = mux_in_sin120;
        10'b0001111001 : logsin2 = mux_in_sin121;
        10'b0001111010 : logsin2 = mux_in_sin122;
        10'b0001111011 : logsin2 = mux_in_sin123;
        10'b0001111100 : logsin2 = mux_in_sin124;
        10'b0001111101 : logsin2 = mux_in_sin125;
        10'b0001111110 : logsin2 = mux_in_sin126;
        10'b0001111111 : logsin2 = mux_in_sin127;
        10'b0010000000 : logsin2 = mux_in_sin128;
        10'b0010000001 : logsin2 = mux_in_sin129;
        10'b0010000010 : logsin2 = mux_in_sin130;
        10'b0010000011 : logsin2 = mux_in_sin131;
        10'b0010000100 : logsin2 = mux_in_sin132;
        10'b0010000101 : logsin2 = mux_in_sin133;
        10'b0010000110 : logsin2 = mux_in_sin134;
        10'b0010000111 : logsin2 = mux_in_sin135;
        10'b0010001000 : logsin2 = mux_in_sin136;
        10'b0010001001 : logsin2 = mux_in_sin137;
        10'b0010001010 : logsin2 = mux_in_sin138;
        10'b0010001011 : logsin2 = mux_in_sin139;
        10'b0010001100 : logsin2 = mux_in_sin140;
        10'b0010001101 : logsin2 = mux_in_sin141;
        10'b0010001110 : logsin2 = mux_in_sin142;
        10'b0010001111 : logsin2 = mux_in_sin143;
        10'b0010010000 : logsin2 = mux_in_sin144;
        10'b0010010001 : logsin2 = mux_in_sin145;
        10'b0010010010 : logsin2 = mux_in_sin146;
        10'b0010010011 : logsin2 = mux_in_sin147;
        10'b0010010100 : logsin2 = mux_in_sin148;
        10'b0010010101 : logsin2 = mux_in_sin149;
        10'b0010010110 : logsin2 = mux_in_sin150;
        10'b0010010111 : logsin2 = mux_in_sin151;
        10'b0010011000 : logsin2 = mux_in_sin152;
        10'b0010011001 : logsin2 = mux_in_sin153;
        10'b0010011010 : logsin2 = mux_in_sin154;
        10'b0010011011 : logsin2 = mux_in_sin155;
        10'b0010011100 : logsin2 = mux_in_sin156;
        10'b0010011101 : logsin2 = mux_in_sin157;
        10'b0010011110 : logsin2 = mux_in_sin158;
        10'b0010011111 : logsin2 = mux_in_sin159;
        10'b0010100000 : logsin2 = mux_in_sin160;
        10'b0010100001 : logsin2 = mux_in_sin161;
        10'b0010100010 : logsin2 = mux_in_sin162;
        10'b0010100011 : logsin2 = mux_in_sin163;
        10'b0010100100 : logsin2 = mux_in_sin164;
        10'b0010100101 : logsin2 = mux_in_sin165;
        10'b0010100110 : logsin2 = mux_in_sin166;
        10'b0010100111 : logsin2 = mux_in_sin167;
        10'b0010101000 : logsin2 = mux_in_sin168;
        10'b0010101001 : logsin2 = mux_in_sin169;
        10'b0010101010 : logsin2 = mux_in_sin170;
        10'b0010101011 : logsin2 = mux_in_sin171;
        10'b0010101100 : logsin2 = mux_in_sin172;
        10'b0010101101 : logsin2 = mux_in_sin173;
        10'b0010101110 : logsin2 = mux_in_sin174;
        10'b0010101111 : logsin2 = mux_in_sin175;
        10'b0010110000 : logsin2 = mux_in_sin176;
        10'b0010110001 : logsin2 = mux_in_sin177;
        10'b0010110010 : logsin2 = mux_in_sin178;
        10'b0010110011 : logsin2 = mux_in_sin179;
        10'b0010110100 : logsin2 = mux_in_sin180;
        10'b0010110101 : logsin2 = mux_in_sin181;
        10'b0010110110 : logsin2 = mux_in_sin182;
        10'b0010110111 : logsin2 = mux_in_sin183;
        10'b0010111000 : logsin2 = mux_in_sin184;
        10'b0010111001 : logsin2 = mux_in_sin185;
        10'b0010111010 : logsin2 = mux_in_sin186;
        10'b0010111011 : logsin2 = mux_in_sin187;
        10'b0010111100 : logsin2 = mux_in_sin188;
        10'b0010111101 : logsin2 = mux_in_sin189;
        10'b0010111110 : logsin2 = mux_in_sin190;
        10'b0010111111 : logsin2 = mux_in_sin191;
        10'b0011000000 : logsin2 = mux_in_sin192;
        10'b0011000001 : logsin2 = mux_in_sin193;
        10'b0011000010 : logsin2 = mux_in_sin194;
        10'b0011000011 : logsin2 = mux_in_sin195;
        10'b0011000100 : logsin2 = mux_in_sin196;
        10'b0011000101 : logsin2 = mux_in_sin197;
        10'b0011000110 : logsin2 = mux_in_sin198;
        10'b0011000111 : logsin2 = mux_in_sin199;
        10'b0011001000 : logsin2 = mux_in_sin200;
        10'b0011001001 : logsin2 = mux_in_sin201;
        10'b0011001010 : logsin2 = mux_in_sin202;
        10'b0011001011 : logsin2 = mux_in_sin203;
        10'b0011001100 : logsin2 = mux_in_sin204;
        10'b0011001101 : logsin2 = mux_in_sin205;
        10'b0011001110 : logsin2 = mux_in_sin206;
        10'b0011001111 : logsin2 = mux_in_sin207;
        10'b0011010000 : logsin2 = mux_in_sin208;
        10'b0011010001 : logsin2 = mux_in_sin209;
        10'b0011010010 : logsin2 = mux_in_sin210;
        10'b0011010011 : logsin2 = mux_in_sin211;
        10'b0011010100 : logsin2 = mux_in_sin212;
        10'b0011010101 : logsin2 = mux_in_sin213;
        10'b0011010110 : logsin2 = mux_in_sin214;
        10'b0011010111 : logsin2 = mux_in_sin215;
        10'b0011011000 : logsin2 = mux_in_sin216;
        10'b0011011001 : logsin2 = mux_in_sin217;
        10'b0011011010 : logsin2 = mux_in_sin218;
        10'b0011011011 : logsin2 = mux_in_sin219;
        10'b0011011100 : logsin2 = mux_in_sin220;
        10'b0011011101 : logsin2 = mux_in_sin221;
        10'b0011011110 : logsin2 = mux_in_sin222;
        10'b0011011111 : logsin2 = mux_in_sin223;
        10'b0011100000 : logsin2 = mux_in_sin224;
        10'b0011100001 : logsin2 = mux_in_sin225;
        10'b0011100010 : logsin2 = mux_in_sin226;
        10'b0011100011 : logsin2 = mux_in_sin227;
        10'b0011100100 : logsin2 = mux_in_sin228;
        10'b0011100101 : logsin2 = mux_in_sin229;
        10'b0011100110 : logsin2 = mux_in_sin230;
        10'b0011100111 : logsin2 = mux_in_sin231;
        10'b0011101000 : logsin2 = mux_in_sin232;
        10'b0011101001 : logsin2 = mux_in_sin233;
        10'b0011101010 : logsin2 = mux_in_sin234;
        10'b0011101011 : logsin2 = mux_in_sin235;
        10'b0011101100 : logsin2 = mux_in_sin236;
        10'b0011101101 : logsin2 = mux_in_sin237;
        10'b0011101110 : logsin2 = mux_in_sin238;
        10'b0011101111 : logsin2 = mux_in_sin239;
        10'b0011110000 : logsin2 = mux_in_sin240;
        10'b0011110001 : logsin2 = mux_in_sin241;
        10'b0011110010 : logsin2 = mux_in_sin242;
        10'b0011110011 : logsin2 = mux_in_sin243;
        10'b0011110100 : logsin2 = mux_in_sin244;
        10'b0011110101 : logsin2 = mux_in_sin245;
        10'b0011110110 : logsin2 = mux_in_sin246;
        10'b0011110111 : logsin2 = mux_in_sin247;
        10'b0011111000 : logsin2 = mux_in_sin248;
        10'b0011111001 : logsin2 = mux_in_sin249;
        10'b0011111010 : logsin2 = mux_in_sin250;
        10'b0011111011 : logsin2 = mux_in_sin251;
        10'b0011111100 : logsin2 = mux_in_sin252;
        10'b0011111101 : logsin2 = mux_in_sin253;
        10'b0011111110 : logsin2 = mux_in_sin254;
        10'b0011111111 : logsin2 = mux_in_sin255;
        10'b0100000000 : logsin2 = mux_in_sin256;
        10'b0100000001 : logsin2 = mux_in_sin257;
        10'b0100000010 : logsin2 = mux_in_sin258;
        10'b0100000011 : logsin2 = mux_in_sin259;
        10'b0100000100 : logsin2 = mux_in_sin260;
        10'b0100000101 : logsin2 = mux_in_sin261;
        10'b0100000110 : logsin2 = mux_in_sin262;
        10'b0100000111 : logsin2 = mux_in_sin263;
        10'b0100001000 : logsin2 = mux_in_sin264;
        10'b0100001001 : logsin2 = mux_in_sin265;
        10'b0100001010 : logsin2 = mux_in_sin266;
        10'b0100001011 : logsin2 = mux_in_sin267;
        10'b0100001100 : logsin2 = mux_in_sin268;
        10'b0100001101 : logsin2 = mux_in_sin269;
        10'b0100001110 : logsin2 = mux_in_sin270;
        10'b0100001111 : logsin2 = mux_in_sin271;
        10'b0100010000 : logsin2 = mux_in_sin272;
        10'b0100010001 : logsin2 = mux_in_sin273;
        10'b0100010010 : logsin2 = mux_in_sin274;
        10'b0100010011 : logsin2 = mux_in_sin275;
        10'b0100010100 : logsin2 = mux_in_sin276;
        10'b0100010101 : logsin2 = mux_in_sin277;
        10'b0100010110 : logsin2 = mux_in_sin278;
        10'b0100010111 : logsin2 = mux_in_sin279;
        10'b0100011000 : logsin2 = mux_in_sin280;
        10'b0100011001 : logsin2 = mux_in_sin281;
        10'b0100011010 : logsin2 = mux_in_sin282;
        10'b0100011011 : logsin2 = mux_in_sin283;
        10'b0100011100 : logsin2 = mux_in_sin284;
        10'b0100011101 : logsin2 = mux_in_sin285;
        10'b0100011110 : logsin2 = mux_in_sin286;
        10'b0100011111 : logsin2 = mux_in_sin287;
        10'b0100100000 : logsin2 = mux_in_sin288;
        10'b0100100001 : logsin2 = mux_in_sin289;
        10'b0100100010 : logsin2 = mux_in_sin290;
        10'b0100100011 : logsin2 = mux_in_sin291;
        10'b0100100100 : logsin2 = mux_in_sin292;
        10'b0100100101 : logsin2 = mux_in_sin293;
        10'b0100100110 : logsin2 = mux_in_sin294;
        10'b0100100111 : logsin2 = mux_in_sin295;
        10'b0100101000 : logsin2 = mux_in_sin296;
        10'b0100101001 : logsin2 = mux_in_sin297;
        10'b0100101010 : logsin2 = mux_in_sin298;
        10'b0100101011 : logsin2 = mux_in_sin299;
        10'b0100101100 : logsin2 = mux_in_sin300;
        10'b0100101101 : logsin2 = mux_in_sin301;
        10'b0100101110 : logsin2 = mux_in_sin302;
        10'b0100101111 : logsin2 = mux_in_sin303;
        10'b0100110000 : logsin2 = mux_in_sin304;
        10'b0100110001 : logsin2 = mux_in_sin305;
        10'b0100110010 : logsin2 = mux_in_sin306;
        10'b0100110011 : logsin2 = mux_in_sin307;
        10'b0100110100 : logsin2 = mux_in_sin308;
        10'b0100110101 : logsin2 = mux_in_sin309;
        10'b0100110110 : logsin2 = mux_in_sin310;
        10'b0100110111 : logsin2 = mux_in_sin311;
        10'b0100111000 : logsin2 = mux_in_sin312;
        10'b0100111001 : logsin2 = mux_in_sin313;
        10'b0100111010 : logsin2 = mux_in_sin314;
        10'b0100111011 : logsin2 = mux_in_sin315;
        10'b0100111100 : logsin2 = mux_in_sin316;
        10'b0100111101 : logsin2 = mux_in_sin317;
        10'b0100111110 : logsin2 = mux_in_sin318;
        10'b0100111111 : logsin2 = mux_in_sin319;
        10'b0101000000 : logsin2 = mux_in_sin320;
        10'b0101000001 : logsin2 = mux_in_sin321;
        10'b0101000010 : logsin2 = mux_in_sin322;
        10'b0101000011 : logsin2 = mux_in_sin323;
        10'b0101000100 : logsin2 = mux_in_sin324;
        10'b0101000101 : logsin2 = mux_in_sin325;
        10'b0101000110 : logsin2 = mux_in_sin326;
        10'b0101000111 : logsin2 = mux_in_sin327;
        10'b0101001000 : logsin2 = mux_in_sin328;
        10'b0101001001 : logsin2 = mux_in_sin329;
        10'b0101001010 : logsin2 = mux_in_sin330;
        10'b0101001011 : logsin2 = mux_in_sin331;
        10'b0101001100 : logsin2 = mux_in_sin332;
        10'b0101001101 : logsin2 = mux_in_sin333;
        10'b0101001110 : logsin2 = mux_in_sin334;
        10'b0101001111 : logsin2 = mux_in_sin335;
        10'b0101010000 : logsin2 = mux_in_sin336;
        10'b0101010001 : logsin2 = mux_in_sin337;
        10'b0101010010 : logsin2 = mux_in_sin338;
        10'b0101010011 : logsin2 = mux_in_sin339;
        10'b0101010100 : logsin2 = mux_in_sin340;
        10'b0101010101 : logsin2 = mux_in_sin341;
        10'b0101010110 : logsin2 = mux_in_sin342;
        10'b0101010111 : logsin2 = mux_in_sin343;
        10'b0101011000 : logsin2 = mux_in_sin344;
        10'b0101011001 : logsin2 = mux_in_sin345;
        10'b0101011010 : logsin2 = mux_in_sin346;
        10'b0101011011 : logsin2 = mux_in_sin347;
        10'b0101011100 : logsin2 = mux_in_sin348;
        10'b0101011101 : logsin2 = mux_in_sin349;
        10'b0101011110 : logsin2 = mux_in_sin350;
        10'b0101011111 : logsin2 = mux_in_sin351;
        10'b0101100000 : logsin2 = mux_in_sin352;
        10'b0101100001 : logsin2 = mux_in_sin353;
        10'b0101100010 : logsin2 = mux_in_sin354;
        10'b0101100011 : logsin2 = mux_in_sin355;
        10'b0101100100 : logsin2 = mux_in_sin356;
        10'b0101100101 : logsin2 = mux_in_sin357;
        10'b0101100110 : logsin2 = mux_in_sin358;
        10'b0101100111 : logsin2 = mux_in_sin359;
        10'b0101101000 : logsin2 = mux_in_sin360;
        10'b0101101001 : logsin2 = mux_in_sin361;
        10'b0101101010 : logsin2 = mux_in_sin362;
        10'b0101101011 : logsin2 = mux_in_sin363;
        10'b0101101100 : logsin2 = mux_in_sin364;
        10'b0101101101 : logsin2 = mux_in_sin365;
        10'b0101101110 : logsin2 = mux_in_sin366;
        10'b0101101111 : logsin2 = mux_in_sin367;
        10'b0101110000 : logsin2 = mux_in_sin368;
        10'b0101110001 : logsin2 = mux_in_sin369;
        10'b0101110010 : logsin2 = mux_in_sin370;
        10'b0101110011 : logsin2 = mux_in_sin371;
        10'b0101110100 : logsin2 = mux_in_sin372;
        10'b0101110101 : logsin2 = mux_in_sin373;
        10'b0101110110 : logsin2 = mux_in_sin374;
        10'b0101110111 : logsin2 = mux_in_sin375;
        10'b0101111000 : logsin2 = mux_in_sin376;
        10'b0101111001 : logsin2 = mux_in_sin377;
        10'b0101111010 : logsin2 = mux_in_sin378;
        10'b0101111011 : logsin2 = mux_in_sin379;
        10'b0101111100 : logsin2 = mux_in_sin380;
        10'b0101111101 : logsin2 = mux_in_sin381;
        10'b0101111110 : logsin2 = mux_in_sin382;
        10'b0101111111 : logsin2 = mux_in_sin383;
        10'b0110000000 : logsin2 = mux_in_sin384;
        10'b0110000001 : logsin2 = mux_in_sin385;
        10'b0110000010 : logsin2 = mux_in_sin386;
        10'b0110000011 : logsin2 = mux_in_sin387;
        10'b0110000100 : logsin2 = mux_in_sin388;
        10'b0110000101 : logsin2 = mux_in_sin389;
        10'b0110000110 : logsin2 = mux_in_sin390;
        10'b0110000111 : logsin2 = mux_in_sin391;
        10'b0110001000 : logsin2 = mux_in_sin392;
        10'b0110001001 : logsin2 = mux_in_sin393;
        10'b0110001010 : logsin2 = mux_in_sin394;
        10'b0110001011 : logsin2 = mux_in_sin395;
        10'b0110001100 : logsin2 = mux_in_sin396;
        10'b0110001101 : logsin2 = mux_in_sin397;
        10'b0110001110 : logsin2 = mux_in_sin398;
        10'b0110001111 : logsin2 = mux_in_sin399;
        10'b0110010000 : logsin2 = mux_in_sin400;
        10'b0110010001 : logsin2 = mux_in_sin401;
        10'b0110010010 : logsin2 = mux_in_sin402;
        10'b0110010011 : logsin2 = mux_in_sin403;
        10'b0110010100 : logsin2 = mux_in_sin404;
        10'b0110010101 : logsin2 = mux_in_sin405;
        10'b0110010110 : logsin2 = mux_in_sin406;
        10'b0110010111 : logsin2 = mux_in_sin407;
        10'b0110011000 : logsin2 = mux_in_sin408;
        10'b0110011001 : logsin2 = mux_in_sin409;
        10'b0110011010 : logsin2 = mux_in_sin410;
        10'b0110011011 : logsin2 = mux_in_sin411;
        10'b0110011100 : logsin2 = mux_in_sin412;
        10'b0110011101 : logsin2 = mux_in_sin413;
        10'b0110011110 : logsin2 = mux_in_sin414;
        10'b0110011111 : logsin2 = mux_in_sin415;
        10'b0110100000 : logsin2 = mux_in_sin416;
        10'b0110100001 : logsin2 = mux_in_sin417;
        10'b0110100010 : logsin2 = mux_in_sin418;
        10'b0110100011 : logsin2 = mux_in_sin419;
        10'b0110100100 : logsin2 = mux_in_sin420;
        10'b0110100101 : logsin2 = mux_in_sin421;
        10'b0110100110 : logsin2 = mux_in_sin422;
        10'b0110100111 : logsin2 = mux_in_sin423;
        10'b0110101000 : logsin2 = mux_in_sin424;
        10'b0110101001 : logsin2 = mux_in_sin425;
        10'b0110101010 : logsin2 = mux_in_sin426;
        10'b0110101011 : logsin2 = mux_in_sin427;
        10'b0110101100 : logsin2 = mux_in_sin428;
        10'b0110101101 : logsin2 = mux_in_sin429;
        10'b0110101110 : logsin2 = mux_in_sin430;
        10'b0110101111 : logsin2 = mux_in_sin431;
        10'b0110110000 : logsin2 = mux_in_sin432;
        10'b0110110001 : logsin2 = mux_in_sin433;
        10'b0110110010 : logsin2 = mux_in_sin434;
        10'b0110110011 : logsin2 = mux_in_sin435;
        10'b0110110100 : logsin2 = mux_in_sin436;
        10'b0110110101 : logsin2 = mux_in_sin437;
        10'b0110110110 : logsin2 = mux_in_sin438;
        10'b0110110111 : logsin2 = mux_in_sin439;
        10'b0110111000 : logsin2 = mux_in_sin440;
        10'b0110111001 : logsin2 = mux_in_sin441;
        10'b0110111010 : logsin2 = mux_in_sin442;
        10'b0110111011 : logsin2 = mux_in_sin443;
        10'b0110111100 : logsin2 = mux_in_sin444;
        10'b0110111101 : logsin2 = mux_in_sin445;
        10'b0110111110 : logsin2 = mux_in_sin446;
        10'b0110111111 : logsin2 = mux_in_sin447;
        10'b0111000000 : logsin2 = mux_in_sin448;
        10'b0111000001 : logsin2 = mux_in_sin449;
        10'b0111000010 : logsin2 = mux_in_sin450;
        10'b0111000011 : logsin2 = mux_in_sin451;
        10'b0111000100 : logsin2 = mux_in_sin452;
        10'b0111000101 : logsin2 = mux_in_sin453;
        10'b0111000110 : logsin2 = mux_in_sin454;
        10'b0111000111 : logsin2 = mux_in_sin455;
        10'b0111001000 : logsin2 = mux_in_sin456;
        10'b0111001001 : logsin2 = mux_in_sin457;
        10'b0111001010 : logsin2 = mux_in_sin458;
        10'b0111001011 : logsin2 = mux_in_sin459;
        10'b0111001100 : logsin2 = mux_in_sin460;
        10'b0111001101 : logsin2 = mux_in_sin461;
        10'b0111001110 : logsin2 = mux_in_sin462;
        10'b0111001111 : logsin2 = mux_in_sin463;
        10'b0111010000 : logsin2 = mux_in_sin464;
        10'b0111010001 : logsin2 = mux_in_sin465;
        10'b0111010010 : logsin2 = mux_in_sin466;
        10'b0111010011 : logsin2 = mux_in_sin467;
        10'b0111010100 : logsin2 = mux_in_sin468;
        10'b0111010101 : logsin2 = mux_in_sin469;
        10'b0111010110 : logsin2 = mux_in_sin470;
        10'b0111010111 : logsin2 = mux_in_sin471;
        10'b0111011000 : logsin2 = mux_in_sin472;
        10'b0111011001 : logsin2 = mux_in_sin473;
        10'b0111011010 : logsin2 = mux_in_sin474;
        10'b0111011011 : logsin2 = mux_in_sin475;
        10'b0111011100 : logsin2 = mux_in_sin476;
        10'b0111011101 : logsin2 = mux_in_sin477;
        10'b0111011110 : logsin2 = mux_in_sin478;
        10'b0111011111 : logsin2 = mux_in_sin479;
        10'b0111100000 : logsin2 = mux_in_sin480;
        10'b0111100001 : logsin2 = mux_in_sin481;
        10'b0111100010 : logsin2 = mux_in_sin482;
        10'b0111100011 : logsin2 = mux_in_sin483;
        10'b0111100100 : logsin2 = mux_in_sin484;
        10'b0111100101 : logsin2 = mux_in_sin485;
        10'b0111100110 : logsin2 = mux_in_sin486;
        10'b0111100111 : logsin2 = mux_in_sin487;
        10'b0111101000 : logsin2 = mux_in_sin488;
        10'b0111101001 : logsin2 = mux_in_sin489;
        10'b0111101010 : logsin2 = mux_in_sin490;
        10'b0111101011 : logsin2 = mux_in_sin491;
        10'b0111101100 : logsin2 = mux_in_sin492;
        10'b0111101101 : logsin2 = mux_in_sin493;
        10'b0111101110 : logsin2 = mux_in_sin494;
        10'b0111101111 : logsin2 = mux_in_sin495;
        10'b0111110000 : logsin2 = mux_in_sin496;
        10'b0111110001 : logsin2 = mux_in_sin497;
        10'b0111110010 : logsin2 = mux_in_sin498;
        10'b0111110011 : logsin2 = mux_in_sin499;
        10'b0111110100 : logsin2 = mux_in_sin500;
        10'b0111110101 : logsin2 = mux_in_sin501;
        10'b0111110110 : logsin2 = mux_in_sin502;
        10'b0111110111 : logsin2 = mux_in_sin503;
        10'b0111111000 : logsin2 = mux_in_sin504;
        10'b0111111001 : logsin2 = mux_in_sin505;
        10'b0111111010 : logsin2 = mux_in_sin506;
        10'b0111111011 : logsin2 = mux_in_sin507;
        10'b0111111100 : logsin2 = mux_in_sin508;
        10'b0111111101 : logsin2 = mux_in_sin509;
        10'b0111111110 : logsin2 = mux_in_sin510;
        10'b0111111111 : logsin2 = mux_in_sin511;
        10'b1000000000 : logsin2 = mux_in_sin512;
        default: logsin2 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in3)
        10'b0000000000 : logsin3 = mux_in_sin0;
        10'b0000000001 : logsin3 = mux_in_sin1;
        10'b0000000010 : logsin3 = mux_in_sin2;
        10'b0000000011 : logsin3 = mux_in_sin3;
        10'b0000000100 : logsin3 = mux_in_sin4;
        10'b0000000101 : logsin3 = mux_in_sin5;
        10'b0000000110 : logsin3 = mux_in_sin6;
        10'b0000000111 : logsin3 = mux_in_sin7;
        10'b0000001000 : logsin3 = mux_in_sin8;
        10'b0000001001 : logsin3 = mux_in_sin9;
        10'b0000001010 : logsin3 = mux_in_sin10;
        10'b0000001011 : logsin3 = mux_in_sin11;
        10'b0000001100 : logsin3 = mux_in_sin12;
        10'b0000001101 : logsin3 = mux_in_sin13;
        10'b0000001110 : logsin3 = mux_in_sin14;
        10'b0000001111 : logsin3 = mux_in_sin15;
        10'b0000010000 : logsin3 = mux_in_sin16;
        10'b0000010001 : logsin3 = mux_in_sin17;
        10'b0000010010 : logsin3 = mux_in_sin18;
        10'b0000010011 : logsin3 = mux_in_sin19;
        10'b0000010100 : logsin3 = mux_in_sin20;
        10'b0000010101 : logsin3 = mux_in_sin21;
        10'b0000010110 : logsin3 = mux_in_sin22;
        10'b0000010111 : logsin3 = mux_in_sin23;
        10'b0000011000 : logsin3 = mux_in_sin24;
        10'b0000011001 : logsin3 = mux_in_sin25;
        10'b0000011010 : logsin3 = mux_in_sin26;
        10'b0000011011 : logsin3 = mux_in_sin27;
        10'b0000011100 : logsin3 = mux_in_sin28;
        10'b0000011101 : logsin3 = mux_in_sin29;
        10'b0000011110 : logsin3 = mux_in_sin30;
        10'b0000011111 : logsin3 = mux_in_sin31;
        10'b0000100000 : logsin3 = mux_in_sin32;
        10'b0000100001 : logsin3 = mux_in_sin33;
        10'b0000100010 : logsin3 = mux_in_sin34;
        10'b0000100011 : logsin3 = mux_in_sin35;
        10'b0000100100 : logsin3 = mux_in_sin36;
        10'b0000100101 : logsin3 = mux_in_sin37;
        10'b0000100110 : logsin3 = mux_in_sin38;
        10'b0000100111 : logsin3 = mux_in_sin39;
        10'b0000101000 : logsin3 = mux_in_sin40;
        10'b0000101001 : logsin3 = mux_in_sin41;
        10'b0000101010 : logsin3 = mux_in_sin42;
        10'b0000101011 : logsin3 = mux_in_sin43;
        10'b0000101100 : logsin3 = mux_in_sin44;
        10'b0000101101 : logsin3 = mux_in_sin45;
        10'b0000101110 : logsin3 = mux_in_sin46;
        10'b0000101111 : logsin3 = mux_in_sin47;
        10'b0000110000 : logsin3 = mux_in_sin48;
        10'b0000110001 : logsin3 = mux_in_sin49;
        10'b0000110010 : logsin3 = mux_in_sin50;
        10'b0000110011 : logsin3 = mux_in_sin51;
        10'b0000110100 : logsin3 = mux_in_sin52;
        10'b0000110101 : logsin3 = mux_in_sin53;
        10'b0000110110 : logsin3 = mux_in_sin54;
        10'b0000110111 : logsin3 = mux_in_sin55;
        10'b0000111000 : logsin3 = mux_in_sin56;
        10'b0000111001 : logsin3 = mux_in_sin57;
        10'b0000111010 : logsin3 = mux_in_sin58;
        10'b0000111011 : logsin3 = mux_in_sin59;
        10'b0000111100 : logsin3 = mux_in_sin60;
        10'b0000111101 : logsin3 = mux_in_sin61;
        10'b0000111110 : logsin3 = mux_in_sin62;
        10'b0000111111 : logsin3 = mux_in_sin63;
        10'b0001000000 : logsin3 = mux_in_sin64;
        10'b0001000001 : logsin3 = mux_in_sin65;
        10'b0001000010 : logsin3 = mux_in_sin66;
        10'b0001000011 : logsin3 = mux_in_sin67;
        10'b0001000100 : logsin3 = mux_in_sin68;
        10'b0001000101 : logsin3 = mux_in_sin69;
        10'b0001000110 : logsin3 = mux_in_sin70;
        10'b0001000111 : logsin3 = mux_in_sin71;
        10'b0001001000 : logsin3 = mux_in_sin72;
        10'b0001001001 : logsin3 = mux_in_sin73;
        10'b0001001010 : logsin3 = mux_in_sin74;
        10'b0001001011 : logsin3 = mux_in_sin75;
        10'b0001001100 : logsin3 = mux_in_sin76;
        10'b0001001101 : logsin3 = mux_in_sin77;
        10'b0001001110 : logsin3 = mux_in_sin78;
        10'b0001001111 : logsin3 = mux_in_sin79;
        10'b0001010000 : logsin3 = mux_in_sin80;
        10'b0001010001 : logsin3 = mux_in_sin81;
        10'b0001010010 : logsin3 = mux_in_sin82;
        10'b0001010011 : logsin3 = mux_in_sin83;
        10'b0001010100 : logsin3 = mux_in_sin84;
        10'b0001010101 : logsin3 = mux_in_sin85;
        10'b0001010110 : logsin3 = mux_in_sin86;
        10'b0001010111 : logsin3 = mux_in_sin87;
        10'b0001011000 : logsin3 = mux_in_sin88;
        10'b0001011001 : logsin3 = mux_in_sin89;
        10'b0001011010 : logsin3 = mux_in_sin90;
        10'b0001011011 : logsin3 = mux_in_sin91;
        10'b0001011100 : logsin3 = mux_in_sin92;
        10'b0001011101 : logsin3 = mux_in_sin93;
        10'b0001011110 : logsin3 = mux_in_sin94;
        10'b0001011111 : logsin3 = mux_in_sin95;
        10'b0001100000 : logsin3 = mux_in_sin96;
        10'b0001100001 : logsin3 = mux_in_sin97;
        10'b0001100010 : logsin3 = mux_in_sin98;
        10'b0001100011 : logsin3 = mux_in_sin99;
        10'b0001100100 : logsin3 = mux_in_sin100;
        10'b0001100101 : logsin3 = mux_in_sin101;
        10'b0001100110 : logsin3 = mux_in_sin102;
        10'b0001100111 : logsin3 = mux_in_sin103;
        10'b0001101000 : logsin3 = mux_in_sin104;
        10'b0001101001 : logsin3 = mux_in_sin105;
        10'b0001101010 : logsin3 = mux_in_sin106;
        10'b0001101011 : logsin3 = mux_in_sin107;
        10'b0001101100 : logsin3 = mux_in_sin108;
        10'b0001101101 : logsin3 = mux_in_sin109;
        10'b0001101110 : logsin3 = mux_in_sin110;
        10'b0001101111 : logsin3 = mux_in_sin111;
        10'b0001110000 : logsin3 = mux_in_sin112;
        10'b0001110001 : logsin3 = mux_in_sin113;
        10'b0001110010 : logsin3 = mux_in_sin114;
        10'b0001110011 : logsin3 = mux_in_sin115;
        10'b0001110100 : logsin3 = mux_in_sin116;
        10'b0001110101 : logsin3 = mux_in_sin117;
        10'b0001110110 : logsin3 = mux_in_sin118;
        10'b0001110111 : logsin3 = mux_in_sin119;
        10'b0001111000 : logsin3 = mux_in_sin120;
        10'b0001111001 : logsin3 = mux_in_sin121;
        10'b0001111010 : logsin3 = mux_in_sin122;
        10'b0001111011 : logsin3 = mux_in_sin123;
        10'b0001111100 : logsin3 = mux_in_sin124;
        10'b0001111101 : logsin3 = mux_in_sin125;
        10'b0001111110 : logsin3 = mux_in_sin126;
        10'b0001111111 : logsin3 = mux_in_sin127;
        10'b0010000000 : logsin3 = mux_in_sin128;
        10'b0010000001 : logsin3 = mux_in_sin129;
        10'b0010000010 : logsin3 = mux_in_sin130;
        10'b0010000011 : logsin3 = mux_in_sin131;
        10'b0010000100 : logsin3 = mux_in_sin132;
        10'b0010000101 : logsin3 = mux_in_sin133;
        10'b0010000110 : logsin3 = mux_in_sin134;
        10'b0010000111 : logsin3 = mux_in_sin135;
        10'b0010001000 : logsin3 = mux_in_sin136;
        10'b0010001001 : logsin3 = mux_in_sin137;
        10'b0010001010 : logsin3 = mux_in_sin138;
        10'b0010001011 : logsin3 = mux_in_sin139;
        10'b0010001100 : logsin3 = mux_in_sin140;
        10'b0010001101 : logsin3 = mux_in_sin141;
        10'b0010001110 : logsin3 = mux_in_sin142;
        10'b0010001111 : logsin3 = mux_in_sin143;
        10'b0010010000 : logsin3 = mux_in_sin144;
        10'b0010010001 : logsin3 = mux_in_sin145;
        10'b0010010010 : logsin3 = mux_in_sin146;
        10'b0010010011 : logsin3 = mux_in_sin147;
        10'b0010010100 : logsin3 = mux_in_sin148;
        10'b0010010101 : logsin3 = mux_in_sin149;
        10'b0010010110 : logsin3 = mux_in_sin150;
        10'b0010010111 : logsin3 = mux_in_sin151;
        10'b0010011000 : logsin3 = mux_in_sin152;
        10'b0010011001 : logsin3 = mux_in_sin153;
        10'b0010011010 : logsin3 = mux_in_sin154;
        10'b0010011011 : logsin3 = mux_in_sin155;
        10'b0010011100 : logsin3 = mux_in_sin156;
        10'b0010011101 : logsin3 = mux_in_sin157;
        10'b0010011110 : logsin3 = mux_in_sin158;
        10'b0010011111 : logsin3 = mux_in_sin159;
        10'b0010100000 : logsin3 = mux_in_sin160;
        10'b0010100001 : logsin3 = mux_in_sin161;
        10'b0010100010 : logsin3 = mux_in_sin162;
        10'b0010100011 : logsin3 = mux_in_sin163;
        10'b0010100100 : logsin3 = mux_in_sin164;
        10'b0010100101 : logsin3 = mux_in_sin165;
        10'b0010100110 : logsin3 = mux_in_sin166;
        10'b0010100111 : logsin3 = mux_in_sin167;
        10'b0010101000 : logsin3 = mux_in_sin168;
        10'b0010101001 : logsin3 = mux_in_sin169;
        10'b0010101010 : logsin3 = mux_in_sin170;
        10'b0010101011 : logsin3 = mux_in_sin171;
        10'b0010101100 : logsin3 = mux_in_sin172;
        10'b0010101101 : logsin3 = mux_in_sin173;
        10'b0010101110 : logsin3 = mux_in_sin174;
        10'b0010101111 : logsin3 = mux_in_sin175;
        10'b0010110000 : logsin3 = mux_in_sin176;
        10'b0010110001 : logsin3 = mux_in_sin177;
        10'b0010110010 : logsin3 = mux_in_sin178;
        10'b0010110011 : logsin3 = mux_in_sin179;
        10'b0010110100 : logsin3 = mux_in_sin180;
        10'b0010110101 : logsin3 = mux_in_sin181;
        10'b0010110110 : logsin3 = mux_in_sin182;
        10'b0010110111 : logsin3 = mux_in_sin183;
        10'b0010111000 : logsin3 = mux_in_sin184;
        10'b0010111001 : logsin3 = mux_in_sin185;
        10'b0010111010 : logsin3 = mux_in_sin186;
        10'b0010111011 : logsin3 = mux_in_sin187;
        10'b0010111100 : logsin3 = mux_in_sin188;
        10'b0010111101 : logsin3 = mux_in_sin189;
        10'b0010111110 : logsin3 = mux_in_sin190;
        10'b0010111111 : logsin3 = mux_in_sin191;
        10'b0011000000 : logsin3 = mux_in_sin192;
        10'b0011000001 : logsin3 = mux_in_sin193;
        10'b0011000010 : logsin3 = mux_in_sin194;
        10'b0011000011 : logsin3 = mux_in_sin195;
        10'b0011000100 : logsin3 = mux_in_sin196;
        10'b0011000101 : logsin3 = mux_in_sin197;
        10'b0011000110 : logsin3 = mux_in_sin198;
        10'b0011000111 : logsin3 = mux_in_sin199;
        10'b0011001000 : logsin3 = mux_in_sin200;
        10'b0011001001 : logsin3 = mux_in_sin201;
        10'b0011001010 : logsin3 = mux_in_sin202;
        10'b0011001011 : logsin3 = mux_in_sin203;
        10'b0011001100 : logsin3 = mux_in_sin204;
        10'b0011001101 : logsin3 = mux_in_sin205;
        10'b0011001110 : logsin3 = mux_in_sin206;
        10'b0011001111 : logsin3 = mux_in_sin207;
        10'b0011010000 : logsin3 = mux_in_sin208;
        10'b0011010001 : logsin3 = mux_in_sin209;
        10'b0011010010 : logsin3 = mux_in_sin210;
        10'b0011010011 : logsin3 = mux_in_sin211;
        10'b0011010100 : logsin3 = mux_in_sin212;
        10'b0011010101 : logsin3 = mux_in_sin213;
        10'b0011010110 : logsin3 = mux_in_sin214;
        10'b0011010111 : logsin3 = mux_in_sin215;
        10'b0011011000 : logsin3 = mux_in_sin216;
        10'b0011011001 : logsin3 = mux_in_sin217;
        10'b0011011010 : logsin3 = mux_in_sin218;
        10'b0011011011 : logsin3 = mux_in_sin219;
        10'b0011011100 : logsin3 = mux_in_sin220;
        10'b0011011101 : logsin3 = mux_in_sin221;
        10'b0011011110 : logsin3 = mux_in_sin222;
        10'b0011011111 : logsin3 = mux_in_sin223;
        10'b0011100000 : logsin3 = mux_in_sin224;
        10'b0011100001 : logsin3 = mux_in_sin225;
        10'b0011100010 : logsin3 = mux_in_sin226;
        10'b0011100011 : logsin3 = mux_in_sin227;
        10'b0011100100 : logsin3 = mux_in_sin228;
        10'b0011100101 : logsin3 = mux_in_sin229;
        10'b0011100110 : logsin3 = mux_in_sin230;
        10'b0011100111 : logsin3 = mux_in_sin231;
        10'b0011101000 : logsin3 = mux_in_sin232;
        10'b0011101001 : logsin3 = mux_in_sin233;
        10'b0011101010 : logsin3 = mux_in_sin234;
        10'b0011101011 : logsin3 = mux_in_sin235;
        10'b0011101100 : logsin3 = mux_in_sin236;
        10'b0011101101 : logsin3 = mux_in_sin237;
        10'b0011101110 : logsin3 = mux_in_sin238;
        10'b0011101111 : logsin3 = mux_in_sin239;
        10'b0011110000 : logsin3 = mux_in_sin240;
        10'b0011110001 : logsin3 = mux_in_sin241;
        10'b0011110010 : logsin3 = mux_in_sin242;
        10'b0011110011 : logsin3 = mux_in_sin243;
        10'b0011110100 : logsin3 = mux_in_sin244;
        10'b0011110101 : logsin3 = mux_in_sin245;
        10'b0011110110 : logsin3 = mux_in_sin246;
        10'b0011110111 : logsin3 = mux_in_sin247;
        10'b0011111000 : logsin3 = mux_in_sin248;
        10'b0011111001 : logsin3 = mux_in_sin249;
        10'b0011111010 : logsin3 = mux_in_sin250;
        10'b0011111011 : logsin3 = mux_in_sin251;
        10'b0011111100 : logsin3 = mux_in_sin252;
        10'b0011111101 : logsin3 = mux_in_sin253;
        10'b0011111110 : logsin3 = mux_in_sin254;
        10'b0011111111 : logsin3 = mux_in_sin255;
        10'b0100000000 : logsin3 = mux_in_sin256;
        10'b0100000001 : logsin3 = mux_in_sin257;
        10'b0100000010 : logsin3 = mux_in_sin258;
        10'b0100000011 : logsin3 = mux_in_sin259;
        10'b0100000100 : logsin3 = mux_in_sin260;
        10'b0100000101 : logsin3 = mux_in_sin261;
        10'b0100000110 : logsin3 = mux_in_sin262;
        10'b0100000111 : logsin3 = mux_in_sin263;
        10'b0100001000 : logsin3 = mux_in_sin264;
        10'b0100001001 : logsin3 = mux_in_sin265;
        10'b0100001010 : logsin3 = mux_in_sin266;
        10'b0100001011 : logsin3 = mux_in_sin267;
        10'b0100001100 : logsin3 = mux_in_sin268;
        10'b0100001101 : logsin3 = mux_in_sin269;
        10'b0100001110 : logsin3 = mux_in_sin270;
        10'b0100001111 : logsin3 = mux_in_sin271;
        10'b0100010000 : logsin3 = mux_in_sin272;
        10'b0100010001 : logsin3 = mux_in_sin273;
        10'b0100010010 : logsin3 = mux_in_sin274;
        10'b0100010011 : logsin3 = mux_in_sin275;
        10'b0100010100 : logsin3 = mux_in_sin276;
        10'b0100010101 : logsin3 = mux_in_sin277;
        10'b0100010110 : logsin3 = mux_in_sin278;
        10'b0100010111 : logsin3 = mux_in_sin279;
        10'b0100011000 : logsin3 = mux_in_sin280;
        10'b0100011001 : logsin3 = mux_in_sin281;
        10'b0100011010 : logsin3 = mux_in_sin282;
        10'b0100011011 : logsin3 = mux_in_sin283;
        10'b0100011100 : logsin3 = mux_in_sin284;
        10'b0100011101 : logsin3 = mux_in_sin285;
        10'b0100011110 : logsin3 = mux_in_sin286;
        10'b0100011111 : logsin3 = mux_in_sin287;
        10'b0100100000 : logsin3 = mux_in_sin288;
        10'b0100100001 : logsin3 = mux_in_sin289;
        10'b0100100010 : logsin3 = mux_in_sin290;
        10'b0100100011 : logsin3 = mux_in_sin291;
        10'b0100100100 : logsin3 = mux_in_sin292;
        10'b0100100101 : logsin3 = mux_in_sin293;
        10'b0100100110 : logsin3 = mux_in_sin294;
        10'b0100100111 : logsin3 = mux_in_sin295;
        10'b0100101000 : logsin3 = mux_in_sin296;
        10'b0100101001 : logsin3 = mux_in_sin297;
        10'b0100101010 : logsin3 = mux_in_sin298;
        10'b0100101011 : logsin3 = mux_in_sin299;
        10'b0100101100 : logsin3 = mux_in_sin300;
        10'b0100101101 : logsin3 = mux_in_sin301;
        10'b0100101110 : logsin3 = mux_in_sin302;
        10'b0100101111 : logsin3 = mux_in_sin303;
        10'b0100110000 : logsin3 = mux_in_sin304;
        10'b0100110001 : logsin3 = mux_in_sin305;
        10'b0100110010 : logsin3 = mux_in_sin306;
        10'b0100110011 : logsin3 = mux_in_sin307;
        10'b0100110100 : logsin3 = mux_in_sin308;
        10'b0100110101 : logsin3 = mux_in_sin309;
        10'b0100110110 : logsin3 = mux_in_sin310;
        10'b0100110111 : logsin3 = mux_in_sin311;
        10'b0100111000 : logsin3 = mux_in_sin312;
        10'b0100111001 : logsin3 = mux_in_sin313;
        10'b0100111010 : logsin3 = mux_in_sin314;
        10'b0100111011 : logsin3 = mux_in_sin315;
        10'b0100111100 : logsin3 = mux_in_sin316;
        10'b0100111101 : logsin3 = mux_in_sin317;
        10'b0100111110 : logsin3 = mux_in_sin318;
        10'b0100111111 : logsin3 = mux_in_sin319;
        10'b0101000000 : logsin3 = mux_in_sin320;
        10'b0101000001 : logsin3 = mux_in_sin321;
        10'b0101000010 : logsin3 = mux_in_sin322;
        10'b0101000011 : logsin3 = mux_in_sin323;
        10'b0101000100 : logsin3 = mux_in_sin324;
        10'b0101000101 : logsin3 = mux_in_sin325;
        10'b0101000110 : logsin3 = mux_in_sin326;
        10'b0101000111 : logsin3 = mux_in_sin327;
        10'b0101001000 : logsin3 = mux_in_sin328;
        10'b0101001001 : logsin3 = mux_in_sin329;
        10'b0101001010 : logsin3 = mux_in_sin330;
        10'b0101001011 : logsin3 = mux_in_sin331;
        10'b0101001100 : logsin3 = mux_in_sin332;
        10'b0101001101 : logsin3 = mux_in_sin333;
        10'b0101001110 : logsin3 = mux_in_sin334;
        10'b0101001111 : logsin3 = mux_in_sin335;
        10'b0101010000 : logsin3 = mux_in_sin336;
        10'b0101010001 : logsin3 = mux_in_sin337;
        10'b0101010010 : logsin3 = mux_in_sin338;
        10'b0101010011 : logsin3 = mux_in_sin339;
        10'b0101010100 : logsin3 = mux_in_sin340;
        10'b0101010101 : logsin3 = mux_in_sin341;
        10'b0101010110 : logsin3 = mux_in_sin342;
        10'b0101010111 : logsin3 = mux_in_sin343;
        10'b0101011000 : logsin3 = mux_in_sin344;
        10'b0101011001 : logsin3 = mux_in_sin345;
        10'b0101011010 : logsin3 = mux_in_sin346;
        10'b0101011011 : logsin3 = mux_in_sin347;
        10'b0101011100 : logsin3 = mux_in_sin348;
        10'b0101011101 : logsin3 = mux_in_sin349;
        10'b0101011110 : logsin3 = mux_in_sin350;
        10'b0101011111 : logsin3 = mux_in_sin351;
        10'b0101100000 : logsin3 = mux_in_sin352;
        10'b0101100001 : logsin3 = mux_in_sin353;
        10'b0101100010 : logsin3 = mux_in_sin354;
        10'b0101100011 : logsin3 = mux_in_sin355;
        10'b0101100100 : logsin3 = mux_in_sin356;
        10'b0101100101 : logsin3 = mux_in_sin357;
        10'b0101100110 : logsin3 = mux_in_sin358;
        10'b0101100111 : logsin3 = mux_in_sin359;
        10'b0101101000 : logsin3 = mux_in_sin360;
        10'b0101101001 : logsin3 = mux_in_sin361;
        10'b0101101010 : logsin3 = mux_in_sin362;
        10'b0101101011 : logsin3 = mux_in_sin363;
        10'b0101101100 : logsin3 = mux_in_sin364;
        10'b0101101101 : logsin3 = mux_in_sin365;
        10'b0101101110 : logsin3 = mux_in_sin366;
        10'b0101101111 : logsin3 = mux_in_sin367;
        10'b0101110000 : logsin3 = mux_in_sin368;
        10'b0101110001 : logsin3 = mux_in_sin369;
        10'b0101110010 : logsin3 = mux_in_sin370;
        10'b0101110011 : logsin3 = mux_in_sin371;
        10'b0101110100 : logsin3 = mux_in_sin372;
        10'b0101110101 : logsin3 = mux_in_sin373;
        10'b0101110110 : logsin3 = mux_in_sin374;
        10'b0101110111 : logsin3 = mux_in_sin375;
        10'b0101111000 : logsin3 = mux_in_sin376;
        10'b0101111001 : logsin3 = mux_in_sin377;
        10'b0101111010 : logsin3 = mux_in_sin378;
        10'b0101111011 : logsin3 = mux_in_sin379;
        10'b0101111100 : logsin3 = mux_in_sin380;
        10'b0101111101 : logsin3 = mux_in_sin381;
        10'b0101111110 : logsin3 = mux_in_sin382;
        10'b0101111111 : logsin3 = mux_in_sin383;
        10'b0110000000 : logsin3 = mux_in_sin384;
        10'b0110000001 : logsin3 = mux_in_sin385;
        10'b0110000010 : logsin3 = mux_in_sin386;
        10'b0110000011 : logsin3 = mux_in_sin387;
        10'b0110000100 : logsin3 = mux_in_sin388;
        10'b0110000101 : logsin3 = mux_in_sin389;
        10'b0110000110 : logsin3 = mux_in_sin390;
        10'b0110000111 : logsin3 = mux_in_sin391;
        10'b0110001000 : logsin3 = mux_in_sin392;
        10'b0110001001 : logsin3 = mux_in_sin393;
        10'b0110001010 : logsin3 = mux_in_sin394;
        10'b0110001011 : logsin3 = mux_in_sin395;
        10'b0110001100 : logsin3 = mux_in_sin396;
        10'b0110001101 : logsin3 = mux_in_sin397;
        10'b0110001110 : logsin3 = mux_in_sin398;
        10'b0110001111 : logsin3 = mux_in_sin399;
        10'b0110010000 : logsin3 = mux_in_sin400;
        10'b0110010001 : logsin3 = mux_in_sin401;
        10'b0110010010 : logsin3 = mux_in_sin402;
        10'b0110010011 : logsin3 = mux_in_sin403;
        10'b0110010100 : logsin3 = mux_in_sin404;
        10'b0110010101 : logsin3 = mux_in_sin405;
        10'b0110010110 : logsin3 = mux_in_sin406;
        10'b0110010111 : logsin3 = mux_in_sin407;
        10'b0110011000 : logsin3 = mux_in_sin408;
        10'b0110011001 : logsin3 = mux_in_sin409;
        10'b0110011010 : logsin3 = mux_in_sin410;
        10'b0110011011 : logsin3 = mux_in_sin411;
        10'b0110011100 : logsin3 = mux_in_sin412;
        10'b0110011101 : logsin3 = mux_in_sin413;
        10'b0110011110 : logsin3 = mux_in_sin414;
        10'b0110011111 : logsin3 = mux_in_sin415;
        10'b0110100000 : logsin3 = mux_in_sin416;
        10'b0110100001 : logsin3 = mux_in_sin417;
        10'b0110100010 : logsin3 = mux_in_sin418;
        10'b0110100011 : logsin3 = mux_in_sin419;
        10'b0110100100 : logsin3 = mux_in_sin420;
        10'b0110100101 : logsin3 = mux_in_sin421;
        10'b0110100110 : logsin3 = mux_in_sin422;
        10'b0110100111 : logsin3 = mux_in_sin423;
        10'b0110101000 : logsin3 = mux_in_sin424;
        10'b0110101001 : logsin3 = mux_in_sin425;
        10'b0110101010 : logsin3 = mux_in_sin426;
        10'b0110101011 : logsin3 = mux_in_sin427;
        10'b0110101100 : logsin3 = mux_in_sin428;
        10'b0110101101 : logsin3 = mux_in_sin429;
        10'b0110101110 : logsin3 = mux_in_sin430;
        10'b0110101111 : logsin3 = mux_in_sin431;
        10'b0110110000 : logsin3 = mux_in_sin432;
        10'b0110110001 : logsin3 = mux_in_sin433;
        10'b0110110010 : logsin3 = mux_in_sin434;
        10'b0110110011 : logsin3 = mux_in_sin435;
        10'b0110110100 : logsin3 = mux_in_sin436;
        10'b0110110101 : logsin3 = mux_in_sin437;
        10'b0110110110 : logsin3 = mux_in_sin438;
        10'b0110110111 : logsin3 = mux_in_sin439;
        10'b0110111000 : logsin3 = mux_in_sin440;
        10'b0110111001 : logsin3 = mux_in_sin441;
        10'b0110111010 : logsin3 = mux_in_sin442;
        10'b0110111011 : logsin3 = mux_in_sin443;
        10'b0110111100 : logsin3 = mux_in_sin444;
        10'b0110111101 : logsin3 = mux_in_sin445;
        10'b0110111110 : logsin3 = mux_in_sin446;
        10'b0110111111 : logsin3 = mux_in_sin447;
        10'b0111000000 : logsin3 = mux_in_sin448;
        10'b0111000001 : logsin3 = mux_in_sin449;
        10'b0111000010 : logsin3 = mux_in_sin450;
        10'b0111000011 : logsin3 = mux_in_sin451;
        10'b0111000100 : logsin3 = mux_in_sin452;
        10'b0111000101 : logsin3 = mux_in_sin453;
        10'b0111000110 : logsin3 = mux_in_sin454;
        10'b0111000111 : logsin3 = mux_in_sin455;
        10'b0111001000 : logsin3 = mux_in_sin456;
        10'b0111001001 : logsin3 = mux_in_sin457;
        10'b0111001010 : logsin3 = mux_in_sin458;
        10'b0111001011 : logsin3 = mux_in_sin459;
        10'b0111001100 : logsin3 = mux_in_sin460;
        10'b0111001101 : logsin3 = mux_in_sin461;
        10'b0111001110 : logsin3 = mux_in_sin462;
        10'b0111001111 : logsin3 = mux_in_sin463;
        10'b0111010000 : logsin3 = mux_in_sin464;
        10'b0111010001 : logsin3 = mux_in_sin465;
        10'b0111010010 : logsin3 = mux_in_sin466;
        10'b0111010011 : logsin3 = mux_in_sin467;
        10'b0111010100 : logsin3 = mux_in_sin468;
        10'b0111010101 : logsin3 = mux_in_sin469;
        10'b0111010110 : logsin3 = mux_in_sin470;
        10'b0111010111 : logsin3 = mux_in_sin471;
        10'b0111011000 : logsin3 = mux_in_sin472;
        10'b0111011001 : logsin3 = mux_in_sin473;
        10'b0111011010 : logsin3 = mux_in_sin474;
        10'b0111011011 : logsin3 = mux_in_sin475;
        10'b0111011100 : logsin3 = mux_in_sin476;
        10'b0111011101 : logsin3 = mux_in_sin477;
        10'b0111011110 : logsin3 = mux_in_sin478;
        10'b0111011111 : logsin3 = mux_in_sin479;
        10'b0111100000 : logsin3 = mux_in_sin480;
        10'b0111100001 : logsin3 = mux_in_sin481;
        10'b0111100010 : logsin3 = mux_in_sin482;
        10'b0111100011 : logsin3 = mux_in_sin483;
        10'b0111100100 : logsin3 = mux_in_sin484;
        10'b0111100101 : logsin3 = mux_in_sin485;
        10'b0111100110 : logsin3 = mux_in_sin486;
        10'b0111100111 : logsin3 = mux_in_sin487;
        10'b0111101000 : logsin3 = mux_in_sin488;
        10'b0111101001 : logsin3 = mux_in_sin489;
        10'b0111101010 : logsin3 = mux_in_sin490;
        10'b0111101011 : logsin3 = mux_in_sin491;
        10'b0111101100 : logsin3 = mux_in_sin492;
        10'b0111101101 : logsin3 = mux_in_sin493;
        10'b0111101110 : logsin3 = mux_in_sin494;
        10'b0111101111 : logsin3 = mux_in_sin495;
        10'b0111110000 : logsin3 = mux_in_sin496;
        10'b0111110001 : logsin3 = mux_in_sin497;
        10'b0111110010 : logsin3 = mux_in_sin498;
        10'b0111110011 : logsin3 = mux_in_sin499;
        10'b0111110100 : logsin3 = mux_in_sin500;
        10'b0111110101 : logsin3 = mux_in_sin501;
        10'b0111110110 : logsin3 = mux_in_sin502;
        10'b0111110111 : logsin3 = mux_in_sin503;
        10'b0111111000 : logsin3 = mux_in_sin504;
        10'b0111111001 : logsin3 = mux_in_sin505;
        10'b0111111010 : logsin3 = mux_in_sin506;
        10'b0111111011 : logsin3 = mux_in_sin507;
        10'b0111111100 : logsin3 = mux_in_sin508;
        10'b0111111101 : logsin3 = mux_in_sin509;
        10'b0111111110 : logsin3 = mux_in_sin510;
        10'b0111111111 : logsin3 = mux_in_sin511;
        10'b1000000000 : logsin3 = mux_in_sin512;
        default: logsin3 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in1)
        10'b0000000000 : logcos1 = mux_in_cos0;
        10'b0000000001 : logcos1 = mux_in_cos1;
        10'b0000000010 : logcos1 = mux_in_cos2;
        10'b0000000011 : logcos1 = mux_in_cos3;
        10'b0000000100 : logcos1 = mux_in_cos4;
        10'b0000000101 : logcos1 = mux_in_cos5;
        10'b0000000110 : logcos1 = mux_in_cos6;
        10'b0000000111 : logcos1 = mux_in_cos7;
        10'b0000001000 : logcos1 = mux_in_cos8;
        10'b0000001001 : logcos1 = mux_in_cos9;
        10'b0000001010 : logcos1 = mux_in_cos10;
        10'b0000001011 : logcos1 = mux_in_cos11;
        10'b0000001100 : logcos1 = mux_in_cos12;
        10'b0000001101 : logcos1 = mux_in_cos13;
        10'b0000001110 : logcos1 = mux_in_cos14;
        10'b0000001111 : logcos1 = mux_in_cos15;
        10'b0000010000 : logcos1 = mux_in_cos16;
        10'b0000010001 : logcos1 = mux_in_cos17;
        10'b0000010010 : logcos1 = mux_in_cos18;
        10'b0000010011 : logcos1 = mux_in_cos19;
        10'b0000010100 : logcos1 = mux_in_cos20;
        10'b0000010101 : logcos1 = mux_in_cos21;
        10'b0000010110 : logcos1 = mux_in_cos22;
        10'b0000010111 : logcos1 = mux_in_cos23;
        10'b0000011000 : logcos1 = mux_in_cos24;
        10'b0000011001 : logcos1 = mux_in_cos25;
        10'b0000011010 : logcos1 = mux_in_cos26;
        10'b0000011011 : logcos1 = mux_in_cos27;
        10'b0000011100 : logcos1 = mux_in_cos28;
        10'b0000011101 : logcos1 = mux_in_cos29;
        10'b0000011110 : logcos1 = mux_in_cos30;
        10'b0000011111 : logcos1 = mux_in_cos31;
        10'b0000100000 : logcos1 = mux_in_cos32;
        10'b0000100001 : logcos1 = mux_in_cos33;
        10'b0000100010 : logcos1 = mux_in_cos34;
        10'b0000100011 : logcos1 = mux_in_cos35;
        10'b0000100100 : logcos1 = mux_in_cos36;
        10'b0000100101 : logcos1 = mux_in_cos37;
        10'b0000100110 : logcos1 = mux_in_cos38;
        10'b0000100111 : logcos1 = mux_in_cos39;
        10'b0000101000 : logcos1 = mux_in_cos40;
        10'b0000101001 : logcos1 = mux_in_cos41;
        10'b0000101010 : logcos1 = mux_in_cos42;
        10'b0000101011 : logcos1 = mux_in_cos43;
        10'b0000101100 : logcos1 = mux_in_cos44;
        10'b0000101101 : logcos1 = mux_in_cos45;
        10'b0000101110 : logcos1 = mux_in_cos46;
        10'b0000101111 : logcos1 = mux_in_cos47;
        10'b0000110000 : logcos1 = mux_in_cos48;
        10'b0000110001 : logcos1 = mux_in_cos49;
        10'b0000110010 : logcos1 = mux_in_cos50;
        10'b0000110011 : logcos1 = mux_in_cos51;
        10'b0000110100 : logcos1 = mux_in_cos52;
        10'b0000110101 : logcos1 = mux_in_cos53;
        10'b0000110110 : logcos1 = mux_in_cos54;
        10'b0000110111 : logcos1 = mux_in_cos55;
        10'b0000111000 : logcos1 = mux_in_cos56;
        10'b0000111001 : logcos1 = mux_in_cos57;
        10'b0000111010 : logcos1 = mux_in_cos58;
        10'b0000111011 : logcos1 = mux_in_cos59;
        10'b0000111100 : logcos1 = mux_in_cos60;
        10'b0000111101 : logcos1 = mux_in_cos61;
        10'b0000111110 : logcos1 = mux_in_cos62;
        10'b0000111111 : logcos1 = mux_in_cos63;
        10'b0001000000 : logcos1 = mux_in_cos64;
        10'b0001000001 : logcos1 = mux_in_cos65;
        10'b0001000010 : logcos1 = mux_in_cos66;
        10'b0001000011 : logcos1 = mux_in_cos67;
        10'b0001000100 : logcos1 = mux_in_cos68;
        10'b0001000101 : logcos1 = mux_in_cos69;
        10'b0001000110 : logcos1 = mux_in_cos70;
        10'b0001000111 : logcos1 = mux_in_cos71;
        10'b0001001000 : logcos1 = mux_in_cos72;
        10'b0001001001 : logcos1 = mux_in_cos73;
        10'b0001001010 : logcos1 = mux_in_cos74;
        10'b0001001011 : logcos1 = mux_in_cos75;
        10'b0001001100 : logcos1 = mux_in_cos76;
        10'b0001001101 : logcos1 = mux_in_cos77;
        10'b0001001110 : logcos1 = mux_in_cos78;
        10'b0001001111 : logcos1 = mux_in_cos79;
        10'b0001010000 : logcos1 = mux_in_cos80;
        10'b0001010001 : logcos1 = mux_in_cos81;
        10'b0001010010 : logcos1 = mux_in_cos82;
        10'b0001010011 : logcos1 = mux_in_cos83;
        10'b0001010100 : logcos1 = mux_in_cos84;
        10'b0001010101 : logcos1 = mux_in_cos85;
        10'b0001010110 : logcos1 = mux_in_cos86;
        10'b0001010111 : logcos1 = mux_in_cos87;
        10'b0001011000 : logcos1 = mux_in_cos88;
        10'b0001011001 : logcos1 = mux_in_cos89;
        10'b0001011010 : logcos1 = mux_in_cos90;
        10'b0001011011 : logcos1 = mux_in_cos91;
        10'b0001011100 : logcos1 = mux_in_cos92;
        10'b0001011101 : logcos1 = mux_in_cos93;
        10'b0001011110 : logcos1 = mux_in_cos94;
        10'b0001011111 : logcos1 = mux_in_cos95;
        10'b0001100000 : logcos1 = mux_in_cos96;
        10'b0001100001 : logcos1 = mux_in_cos97;
        10'b0001100010 : logcos1 = mux_in_cos98;
        10'b0001100011 : logcos1 = mux_in_cos99;
        10'b0001100100 : logcos1 = mux_in_cos100;
        10'b0001100101 : logcos1 = mux_in_cos101;
        10'b0001100110 : logcos1 = mux_in_cos102;
        10'b0001100111 : logcos1 = mux_in_cos103;
        10'b0001101000 : logcos1 = mux_in_cos104;
        10'b0001101001 : logcos1 = mux_in_cos105;
        10'b0001101010 : logcos1 = mux_in_cos106;
        10'b0001101011 : logcos1 = mux_in_cos107;
        10'b0001101100 : logcos1 = mux_in_cos108;
        10'b0001101101 : logcos1 = mux_in_cos109;
        10'b0001101110 : logcos1 = mux_in_cos110;
        10'b0001101111 : logcos1 = mux_in_cos111;
        10'b0001110000 : logcos1 = mux_in_cos112;
        10'b0001110001 : logcos1 = mux_in_cos113;
        10'b0001110010 : logcos1 = mux_in_cos114;
        10'b0001110011 : logcos1 = mux_in_cos115;
        10'b0001110100 : logcos1 = mux_in_cos116;
        10'b0001110101 : logcos1 = mux_in_cos117;
        10'b0001110110 : logcos1 = mux_in_cos118;
        10'b0001110111 : logcos1 = mux_in_cos119;
        10'b0001111000 : logcos1 = mux_in_cos120;
        10'b0001111001 : logcos1 = mux_in_cos121;
        10'b0001111010 : logcos1 = mux_in_cos122;
        10'b0001111011 : logcos1 = mux_in_cos123;
        10'b0001111100 : logcos1 = mux_in_cos124;
        10'b0001111101 : logcos1 = mux_in_cos125;
        10'b0001111110 : logcos1 = mux_in_cos126;
        10'b0001111111 : logcos1 = mux_in_cos127;
        10'b0010000000 : logcos1 = mux_in_cos128;
        10'b0010000001 : logcos1 = mux_in_cos129;
        10'b0010000010 : logcos1 = mux_in_cos130;
        10'b0010000011 : logcos1 = mux_in_cos131;
        10'b0010000100 : logcos1 = mux_in_cos132;
        10'b0010000101 : logcos1 = mux_in_cos133;
        10'b0010000110 : logcos1 = mux_in_cos134;
        10'b0010000111 : logcos1 = mux_in_cos135;
        10'b0010001000 : logcos1 = mux_in_cos136;
        10'b0010001001 : logcos1 = mux_in_cos137;
        10'b0010001010 : logcos1 = mux_in_cos138;
        10'b0010001011 : logcos1 = mux_in_cos139;
        10'b0010001100 : logcos1 = mux_in_cos140;
        10'b0010001101 : logcos1 = mux_in_cos141;
        10'b0010001110 : logcos1 = mux_in_cos142;
        10'b0010001111 : logcos1 = mux_in_cos143;
        10'b0010010000 : logcos1 = mux_in_cos144;
        10'b0010010001 : logcos1 = mux_in_cos145;
        10'b0010010010 : logcos1 = mux_in_cos146;
        10'b0010010011 : logcos1 = mux_in_cos147;
        10'b0010010100 : logcos1 = mux_in_cos148;
        10'b0010010101 : logcos1 = mux_in_cos149;
        10'b0010010110 : logcos1 = mux_in_cos150;
        10'b0010010111 : logcos1 = mux_in_cos151;
        10'b0010011000 : logcos1 = mux_in_cos152;
        10'b0010011001 : logcos1 = mux_in_cos153;
        10'b0010011010 : logcos1 = mux_in_cos154;
        10'b0010011011 : logcos1 = mux_in_cos155;
        10'b0010011100 : logcos1 = mux_in_cos156;
        10'b0010011101 : logcos1 = mux_in_cos157;
        10'b0010011110 : logcos1 = mux_in_cos158;
        10'b0010011111 : logcos1 = mux_in_cos159;
        10'b0010100000 : logcos1 = mux_in_cos160;
        10'b0010100001 : logcos1 = mux_in_cos161;
        10'b0010100010 : logcos1 = mux_in_cos162;
        10'b0010100011 : logcos1 = mux_in_cos163;
        10'b0010100100 : logcos1 = mux_in_cos164;
        10'b0010100101 : logcos1 = mux_in_cos165;
        10'b0010100110 : logcos1 = mux_in_cos166;
        10'b0010100111 : logcos1 = mux_in_cos167;
        10'b0010101000 : logcos1 = mux_in_cos168;
        10'b0010101001 : logcos1 = mux_in_cos169;
        10'b0010101010 : logcos1 = mux_in_cos170;
        10'b0010101011 : logcos1 = mux_in_cos171;
        10'b0010101100 : logcos1 = mux_in_cos172;
        10'b0010101101 : logcos1 = mux_in_cos173;
        10'b0010101110 : logcos1 = mux_in_cos174;
        10'b0010101111 : logcos1 = mux_in_cos175;
        10'b0010110000 : logcos1 = mux_in_cos176;
        10'b0010110001 : logcos1 = mux_in_cos177;
        10'b0010110010 : logcos1 = mux_in_cos178;
        10'b0010110011 : logcos1 = mux_in_cos179;
        10'b0010110100 : logcos1 = mux_in_cos180;
        10'b0010110101 : logcos1 = mux_in_cos181;
        10'b0010110110 : logcos1 = mux_in_cos182;
        10'b0010110111 : logcos1 = mux_in_cos183;
        10'b0010111000 : logcos1 = mux_in_cos184;
        10'b0010111001 : logcos1 = mux_in_cos185;
        10'b0010111010 : logcos1 = mux_in_cos186;
        10'b0010111011 : logcos1 = mux_in_cos187;
        10'b0010111100 : logcos1 = mux_in_cos188;
        10'b0010111101 : logcos1 = mux_in_cos189;
        10'b0010111110 : logcos1 = mux_in_cos190;
        10'b0010111111 : logcos1 = mux_in_cos191;
        10'b0011000000 : logcos1 = mux_in_cos192;
        10'b0011000001 : logcos1 = mux_in_cos193;
        10'b0011000010 : logcos1 = mux_in_cos194;
        10'b0011000011 : logcos1 = mux_in_cos195;
        10'b0011000100 : logcos1 = mux_in_cos196;
        10'b0011000101 : logcos1 = mux_in_cos197;
        10'b0011000110 : logcos1 = mux_in_cos198;
        10'b0011000111 : logcos1 = mux_in_cos199;
        10'b0011001000 : logcos1 = mux_in_cos200;
        10'b0011001001 : logcos1 = mux_in_cos201;
        10'b0011001010 : logcos1 = mux_in_cos202;
        10'b0011001011 : logcos1 = mux_in_cos203;
        10'b0011001100 : logcos1 = mux_in_cos204;
        10'b0011001101 : logcos1 = mux_in_cos205;
        10'b0011001110 : logcos1 = mux_in_cos206;
        10'b0011001111 : logcos1 = mux_in_cos207;
        10'b0011010000 : logcos1 = mux_in_cos208;
        10'b0011010001 : logcos1 = mux_in_cos209;
        10'b0011010010 : logcos1 = mux_in_cos210;
        10'b0011010011 : logcos1 = mux_in_cos211;
        10'b0011010100 : logcos1 = mux_in_cos212;
        10'b0011010101 : logcos1 = mux_in_cos213;
        10'b0011010110 : logcos1 = mux_in_cos214;
        10'b0011010111 : logcos1 = mux_in_cos215;
        10'b0011011000 : logcos1 = mux_in_cos216;
        10'b0011011001 : logcos1 = mux_in_cos217;
        10'b0011011010 : logcos1 = mux_in_cos218;
        10'b0011011011 : logcos1 = mux_in_cos219;
        10'b0011011100 : logcos1 = mux_in_cos220;
        10'b0011011101 : logcos1 = mux_in_cos221;
        10'b0011011110 : logcos1 = mux_in_cos222;
        10'b0011011111 : logcos1 = mux_in_cos223;
        10'b0011100000 : logcos1 = mux_in_cos224;
        10'b0011100001 : logcos1 = mux_in_cos225;
        10'b0011100010 : logcos1 = mux_in_cos226;
        10'b0011100011 : logcos1 = mux_in_cos227;
        10'b0011100100 : logcos1 = mux_in_cos228;
        10'b0011100101 : logcos1 = mux_in_cos229;
        10'b0011100110 : logcos1 = mux_in_cos230;
        10'b0011100111 : logcos1 = mux_in_cos231;
        10'b0011101000 : logcos1 = mux_in_cos232;
        10'b0011101001 : logcos1 = mux_in_cos233;
        10'b0011101010 : logcos1 = mux_in_cos234;
        10'b0011101011 : logcos1 = mux_in_cos235;
        10'b0011101100 : logcos1 = mux_in_cos236;
        10'b0011101101 : logcos1 = mux_in_cos237;
        10'b0011101110 : logcos1 = mux_in_cos238;
        10'b0011101111 : logcos1 = mux_in_cos239;
        10'b0011110000 : logcos1 = mux_in_cos240;
        10'b0011110001 : logcos1 = mux_in_cos241;
        10'b0011110010 : logcos1 = mux_in_cos242;
        10'b0011110011 : logcos1 = mux_in_cos243;
        10'b0011110100 : logcos1 = mux_in_cos244;
        10'b0011110101 : logcos1 = mux_in_cos245;
        10'b0011110110 : logcos1 = mux_in_cos246;
        10'b0011110111 : logcos1 = mux_in_cos247;
        10'b0011111000 : logcos1 = mux_in_cos248;
        10'b0011111001 : logcos1 = mux_in_cos249;
        10'b0011111010 : logcos1 = mux_in_cos250;
        10'b0011111011 : logcos1 = mux_in_cos251;
        10'b0011111100 : logcos1 = mux_in_cos252;
        10'b0011111101 : logcos1 = mux_in_cos253;
        10'b0011111110 : logcos1 = mux_in_cos254;
        10'b0011111111 : logcos1 = mux_in_cos255;
        10'b0100000000 : logcos1 = mux_in_cos256;
        10'b0100000001 : logcos1 = mux_in_cos257;
        10'b0100000010 : logcos1 = mux_in_cos258;
        10'b0100000011 : logcos1 = mux_in_cos259;
        10'b0100000100 : logcos1 = mux_in_cos260;
        10'b0100000101 : logcos1 = mux_in_cos261;
        10'b0100000110 : logcos1 = mux_in_cos262;
        10'b0100000111 : logcos1 = mux_in_cos263;
        10'b0100001000 : logcos1 = mux_in_cos264;
        10'b0100001001 : logcos1 = mux_in_cos265;
        10'b0100001010 : logcos1 = mux_in_cos266;
        10'b0100001011 : logcos1 = mux_in_cos267;
        10'b0100001100 : logcos1 = mux_in_cos268;
        10'b0100001101 : logcos1 = mux_in_cos269;
        10'b0100001110 : logcos1 = mux_in_cos270;
        10'b0100001111 : logcos1 = mux_in_cos271;
        10'b0100010000 : logcos1 = mux_in_cos272;
        10'b0100010001 : logcos1 = mux_in_cos273;
        10'b0100010010 : logcos1 = mux_in_cos274;
        10'b0100010011 : logcos1 = mux_in_cos275;
        10'b0100010100 : logcos1 = mux_in_cos276;
        10'b0100010101 : logcos1 = mux_in_cos277;
        10'b0100010110 : logcos1 = mux_in_cos278;
        10'b0100010111 : logcos1 = mux_in_cos279;
        10'b0100011000 : logcos1 = mux_in_cos280;
        10'b0100011001 : logcos1 = mux_in_cos281;
        10'b0100011010 : logcos1 = mux_in_cos282;
        10'b0100011011 : logcos1 = mux_in_cos283;
        10'b0100011100 : logcos1 = mux_in_cos284;
        10'b0100011101 : logcos1 = mux_in_cos285;
        10'b0100011110 : logcos1 = mux_in_cos286;
        10'b0100011111 : logcos1 = mux_in_cos287;
        10'b0100100000 : logcos1 = mux_in_cos288;
        10'b0100100001 : logcos1 = mux_in_cos289;
        10'b0100100010 : logcos1 = mux_in_cos290;
        10'b0100100011 : logcos1 = mux_in_cos291;
        10'b0100100100 : logcos1 = mux_in_cos292;
        10'b0100100101 : logcos1 = mux_in_cos293;
        10'b0100100110 : logcos1 = mux_in_cos294;
        10'b0100100111 : logcos1 = mux_in_cos295;
        10'b0100101000 : logcos1 = mux_in_cos296;
        10'b0100101001 : logcos1 = mux_in_cos297;
        10'b0100101010 : logcos1 = mux_in_cos298;
        10'b0100101011 : logcos1 = mux_in_cos299;
        10'b0100101100 : logcos1 = mux_in_cos300;
        10'b0100101101 : logcos1 = mux_in_cos301;
        10'b0100101110 : logcos1 = mux_in_cos302;
        10'b0100101111 : logcos1 = mux_in_cos303;
        10'b0100110000 : logcos1 = mux_in_cos304;
        10'b0100110001 : logcos1 = mux_in_cos305;
        10'b0100110010 : logcos1 = mux_in_cos306;
        10'b0100110011 : logcos1 = mux_in_cos307;
        10'b0100110100 : logcos1 = mux_in_cos308;
        10'b0100110101 : logcos1 = mux_in_cos309;
        10'b0100110110 : logcos1 = mux_in_cos310;
        10'b0100110111 : logcos1 = mux_in_cos311;
        10'b0100111000 : logcos1 = mux_in_cos312;
        10'b0100111001 : logcos1 = mux_in_cos313;
        10'b0100111010 : logcos1 = mux_in_cos314;
        10'b0100111011 : logcos1 = mux_in_cos315;
        10'b0100111100 : logcos1 = mux_in_cos316;
        10'b0100111101 : logcos1 = mux_in_cos317;
        10'b0100111110 : logcos1 = mux_in_cos318;
        10'b0100111111 : logcos1 = mux_in_cos319;
        10'b0101000000 : logcos1 = mux_in_cos320;
        10'b0101000001 : logcos1 = mux_in_cos321;
        10'b0101000010 : logcos1 = mux_in_cos322;
        10'b0101000011 : logcos1 = mux_in_cos323;
        10'b0101000100 : logcos1 = mux_in_cos324;
        10'b0101000101 : logcos1 = mux_in_cos325;
        10'b0101000110 : logcos1 = mux_in_cos326;
        10'b0101000111 : logcos1 = mux_in_cos327;
        10'b0101001000 : logcos1 = mux_in_cos328;
        10'b0101001001 : logcos1 = mux_in_cos329;
        10'b0101001010 : logcos1 = mux_in_cos330;
        10'b0101001011 : logcos1 = mux_in_cos331;
        10'b0101001100 : logcos1 = mux_in_cos332;
        10'b0101001101 : logcos1 = mux_in_cos333;
        10'b0101001110 : logcos1 = mux_in_cos334;
        10'b0101001111 : logcos1 = mux_in_cos335;
        10'b0101010000 : logcos1 = mux_in_cos336;
        10'b0101010001 : logcos1 = mux_in_cos337;
        10'b0101010010 : logcos1 = mux_in_cos338;
        10'b0101010011 : logcos1 = mux_in_cos339;
        10'b0101010100 : logcos1 = mux_in_cos340;
        10'b0101010101 : logcos1 = mux_in_cos341;
        10'b0101010110 : logcos1 = mux_in_cos342;
        10'b0101010111 : logcos1 = mux_in_cos343;
        10'b0101011000 : logcos1 = mux_in_cos344;
        10'b0101011001 : logcos1 = mux_in_cos345;
        10'b0101011010 : logcos1 = mux_in_cos346;
        10'b0101011011 : logcos1 = mux_in_cos347;
        10'b0101011100 : logcos1 = mux_in_cos348;
        10'b0101011101 : logcos1 = mux_in_cos349;
        10'b0101011110 : logcos1 = mux_in_cos350;
        10'b0101011111 : logcos1 = mux_in_cos351;
        10'b0101100000 : logcos1 = mux_in_cos352;
        10'b0101100001 : logcos1 = mux_in_cos353;
        10'b0101100010 : logcos1 = mux_in_cos354;
        10'b0101100011 : logcos1 = mux_in_cos355;
        10'b0101100100 : logcos1 = mux_in_cos356;
        10'b0101100101 : logcos1 = mux_in_cos357;
        10'b0101100110 : logcos1 = mux_in_cos358;
        10'b0101100111 : logcos1 = mux_in_cos359;
        10'b0101101000 : logcos1 = mux_in_cos360;
        10'b0101101001 : logcos1 = mux_in_cos361;
        10'b0101101010 : logcos1 = mux_in_cos362;
        10'b0101101011 : logcos1 = mux_in_cos363;
        10'b0101101100 : logcos1 = mux_in_cos364;
        10'b0101101101 : logcos1 = mux_in_cos365;
        10'b0101101110 : logcos1 = mux_in_cos366;
        10'b0101101111 : logcos1 = mux_in_cos367;
        10'b0101110000 : logcos1 = mux_in_cos368;
        10'b0101110001 : logcos1 = mux_in_cos369;
        10'b0101110010 : logcos1 = mux_in_cos370;
        10'b0101110011 : logcos1 = mux_in_cos371;
        10'b0101110100 : logcos1 = mux_in_cos372;
        10'b0101110101 : logcos1 = mux_in_cos373;
        10'b0101110110 : logcos1 = mux_in_cos374;
        10'b0101110111 : logcos1 = mux_in_cos375;
        10'b0101111000 : logcos1 = mux_in_cos376;
        10'b0101111001 : logcos1 = mux_in_cos377;
        10'b0101111010 : logcos1 = mux_in_cos378;
        10'b0101111011 : logcos1 = mux_in_cos379;
        10'b0101111100 : logcos1 = mux_in_cos380;
        10'b0101111101 : logcos1 = mux_in_cos381;
        10'b0101111110 : logcos1 = mux_in_cos382;
        10'b0101111111 : logcos1 = mux_in_cos383;
        10'b0110000000 : logcos1 = mux_in_cos384;
        10'b0110000001 : logcos1 = mux_in_cos385;
        10'b0110000010 : logcos1 = mux_in_cos386;
        10'b0110000011 : logcos1 = mux_in_cos387;
        10'b0110000100 : logcos1 = mux_in_cos388;
        10'b0110000101 : logcos1 = mux_in_cos389;
        10'b0110000110 : logcos1 = mux_in_cos390;
        10'b0110000111 : logcos1 = mux_in_cos391;
        10'b0110001000 : logcos1 = mux_in_cos392;
        10'b0110001001 : logcos1 = mux_in_cos393;
        10'b0110001010 : logcos1 = mux_in_cos394;
        10'b0110001011 : logcos1 = mux_in_cos395;
        10'b0110001100 : logcos1 = mux_in_cos396;
        10'b0110001101 : logcos1 = mux_in_cos397;
        10'b0110001110 : logcos1 = mux_in_cos398;
        10'b0110001111 : logcos1 = mux_in_cos399;
        10'b0110010000 : logcos1 = mux_in_cos400;
        10'b0110010001 : logcos1 = mux_in_cos401;
        10'b0110010010 : logcos1 = mux_in_cos402;
        10'b0110010011 : logcos1 = mux_in_cos403;
        10'b0110010100 : logcos1 = mux_in_cos404;
        10'b0110010101 : logcos1 = mux_in_cos405;
        10'b0110010110 : logcos1 = mux_in_cos406;
        10'b0110010111 : logcos1 = mux_in_cos407;
        10'b0110011000 : logcos1 = mux_in_cos408;
        10'b0110011001 : logcos1 = mux_in_cos409;
        10'b0110011010 : logcos1 = mux_in_cos410;
        10'b0110011011 : logcos1 = mux_in_cos411;
        10'b0110011100 : logcos1 = mux_in_cos412;
        10'b0110011101 : logcos1 = mux_in_cos413;
        10'b0110011110 : logcos1 = mux_in_cos414;
        10'b0110011111 : logcos1 = mux_in_cos415;
        10'b0110100000 : logcos1 = mux_in_cos416;
        10'b0110100001 : logcos1 = mux_in_cos417;
        10'b0110100010 : logcos1 = mux_in_cos418;
        10'b0110100011 : logcos1 = mux_in_cos419;
        10'b0110100100 : logcos1 = mux_in_cos420;
        10'b0110100101 : logcos1 = mux_in_cos421;
        10'b0110100110 : logcos1 = mux_in_cos422;
        10'b0110100111 : logcos1 = mux_in_cos423;
        10'b0110101000 : logcos1 = mux_in_cos424;
        10'b0110101001 : logcos1 = mux_in_cos425;
        10'b0110101010 : logcos1 = mux_in_cos426;
        10'b0110101011 : logcos1 = mux_in_cos427;
        10'b0110101100 : logcos1 = mux_in_cos428;
        10'b0110101101 : logcos1 = mux_in_cos429;
        10'b0110101110 : logcos1 = mux_in_cos430;
        10'b0110101111 : logcos1 = mux_in_cos431;
        10'b0110110000 : logcos1 = mux_in_cos432;
        10'b0110110001 : logcos1 = mux_in_cos433;
        10'b0110110010 : logcos1 = mux_in_cos434;
        10'b0110110011 : logcos1 = mux_in_cos435;
        10'b0110110100 : logcos1 = mux_in_cos436;
        10'b0110110101 : logcos1 = mux_in_cos437;
        10'b0110110110 : logcos1 = mux_in_cos438;
        10'b0110110111 : logcos1 = mux_in_cos439;
        10'b0110111000 : logcos1 = mux_in_cos440;
        10'b0110111001 : logcos1 = mux_in_cos441;
        10'b0110111010 : logcos1 = mux_in_cos442;
        10'b0110111011 : logcos1 = mux_in_cos443;
        10'b0110111100 : logcos1 = mux_in_cos444;
        10'b0110111101 : logcos1 = mux_in_cos445;
        10'b0110111110 : logcos1 = mux_in_cos446;
        10'b0110111111 : logcos1 = mux_in_cos447;
        10'b0111000000 : logcos1 = mux_in_cos448;
        10'b0111000001 : logcos1 = mux_in_cos449;
        10'b0111000010 : logcos1 = mux_in_cos450;
        10'b0111000011 : logcos1 = mux_in_cos451;
        10'b0111000100 : logcos1 = mux_in_cos452;
        10'b0111000101 : logcos1 = mux_in_cos453;
        10'b0111000110 : logcos1 = mux_in_cos454;
        10'b0111000111 : logcos1 = mux_in_cos455;
        10'b0111001000 : logcos1 = mux_in_cos456;
        10'b0111001001 : logcos1 = mux_in_cos457;
        10'b0111001010 : logcos1 = mux_in_cos458;
        10'b0111001011 : logcos1 = mux_in_cos459;
        10'b0111001100 : logcos1 = mux_in_cos460;
        10'b0111001101 : logcos1 = mux_in_cos461;
        10'b0111001110 : logcos1 = mux_in_cos462;
        10'b0111001111 : logcos1 = mux_in_cos463;
        10'b0111010000 : logcos1 = mux_in_cos464;
        10'b0111010001 : logcos1 = mux_in_cos465;
        10'b0111010010 : logcos1 = mux_in_cos466;
        10'b0111010011 : logcos1 = mux_in_cos467;
        10'b0111010100 : logcos1 = mux_in_cos468;
        10'b0111010101 : logcos1 = mux_in_cos469;
        10'b0111010110 : logcos1 = mux_in_cos470;
        10'b0111010111 : logcos1 = mux_in_cos471;
        10'b0111011000 : logcos1 = mux_in_cos472;
        10'b0111011001 : logcos1 = mux_in_cos473;
        10'b0111011010 : logcos1 = mux_in_cos474;
        10'b0111011011 : logcos1 = mux_in_cos475;
        10'b0111011100 : logcos1 = mux_in_cos476;
        10'b0111011101 : logcos1 = mux_in_cos477;
        10'b0111011110 : logcos1 = mux_in_cos478;
        10'b0111011111 : logcos1 = mux_in_cos479;
        10'b0111100000 : logcos1 = mux_in_cos480;
        10'b0111100001 : logcos1 = mux_in_cos481;
        10'b0111100010 : logcos1 = mux_in_cos482;
        10'b0111100011 : logcos1 = mux_in_cos483;
        10'b0111100100 : logcos1 = mux_in_cos484;
        10'b0111100101 : logcos1 = mux_in_cos485;
        10'b0111100110 : logcos1 = mux_in_cos486;
        10'b0111100111 : logcos1 = mux_in_cos487;
        10'b0111101000 : logcos1 = mux_in_cos488;
        10'b0111101001 : logcos1 = mux_in_cos489;
        10'b0111101010 : logcos1 = mux_in_cos490;
        10'b0111101011 : logcos1 = mux_in_cos491;
        10'b0111101100 : logcos1 = mux_in_cos492;
        10'b0111101101 : logcos1 = mux_in_cos493;
        10'b0111101110 : logcos1 = mux_in_cos494;
        10'b0111101111 : logcos1 = mux_in_cos495;
        10'b0111110000 : logcos1 = mux_in_cos496;
        10'b0111110001 : logcos1 = mux_in_cos497;
        10'b0111110010 : logcos1 = mux_in_cos498;
        10'b0111110011 : logcos1 = mux_in_cos499;
        10'b0111110100 : logcos1 = mux_in_cos500;
        10'b0111110101 : logcos1 = mux_in_cos501;
        10'b0111110110 : logcos1 = mux_in_cos502;
        10'b0111110111 : logcos1 = mux_in_cos503;
        10'b0111111000 : logcos1 = mux_in_cos504;
        10'b0111111001 : logcos1 = mux_in_cos505;
        10'b0111111010 : logcos1 = mux_in_cos506;
        10'b0111111011 : logcos1 = mux_in_cos507;
        10'b0111111100 : logcos1 = mux_in_cos508;
        10'b0111111101 : logcos1 = mux_in_cos509;
        10'b0111111110 : logcos1 = mux_in_cos510;
        10'b0111111111 : logcos1 = mux_in_cos511;
        10'b1000000000 : logcos1 = mux_in_cos512;
        default: logcos1 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in2)
        10'b0000000000 : logcos2 = mux_in_cos0;
        10'b0000000001 : logcos2 = mux_in_cos1;
        10'b0000000010 : logcos2 = mux_in_cos2;
        10'b0000000011 : logcos2 = mux_in_cos3;
        10'b0000000100 : logcos2 = mux_in_cos4;
        10'b0000000101 : logcos2 = mux_in_cos5;
        10'b0000000110 : logcos2 = mux_in_cos6;
        10'b0000000111 : logcos2 = mux_in_cos7;
        10'b0000001000 : logcos2 = mux_in_cos8;
        10'b0000001001 : logcos2 = mux_in_cos9;
        10'b0000001010 : logcos2 = mux_in_cos10;
        10'b0000001011 : logcos2 = mux_in_cos11;
        10'b0000001100 : logcos2 = mux_in_cos12;
        10'b0000001101 : logcos2 = mux_in_cos13;
        10'b0000001110 : logcos2 = mux_in_cos14;
        10'b0000001111 : logcos2 = mux_in_cos15;
        10'b0000010000 : logcos2 = mux_in_cos16;
        10'b0000010001 : logcos2 = mux_in_cos17;
        10'b0000010010 : logcos2 = mux_in_cos18;
        10'b0000010011 : logcos2 = mux_in_cos19;
        10'b0000010100 : logcos2 = mux_in_cos20;
        10'b0000010101 : logcos2 = mux_in_cos21;
        10'b0000010110 : logcos2 = mux_in_cos22;
        10'b0000010111 : logcos2 = mux_in_cos23;
        10'b0000011000 : logcos2 = mux_in_cos24;
        10'b0000011001 : logcos2 = mux_in_cos25;
        10'b0000011010 : logcos2 = mux_in_cos26;
        10'b0000011011 : logcos2 = mux_in_cos27;
        10'b0000011100 : logcos2 = mux_in_cos28;
        10'b0000011101 : logcos2 = mux_in_cos29;
        10'b0000011110 : logcos2 = mux_in_cos30;
        10'b0000011111 : logcos2 = mux_in_cos31;
        10'b0000100000 : logcos2 = mux_in_cos32;
        10'b0000100001 : logcos2 = mux_in_cos33;
        10'b0000100010 : logcos2 = mux_in_cos34;
        10'b0000100011 : logcos2 = mux_in_cos35;
        10'b0000100100 : logcos2 = mux_in_cos36;
        10'b0000100101 : logcos2 = mux_in_cos37;
        10'b0000100110 : logcos2 = mux_in_cos38;
        10'b0000100111 : logcos2 = mux_in_cos39;
        10'b0000101000 : logcos2 = mux_in_cos40;
        10'b0000101001 : logcos2 = mux_in_cos41;
        10'b0000101010 : logcos2 = mux_in_cos42;
        10'b0000101011 : logcos2 = mux_in_cos43;
        10'b0000101100 : logcos2 = mux_in_cos44;
        10'b0000101101 : logcos2 = mux_in_cos45;
        10'b0000101110 : logcos2 = mux_in_cos46;
        10'b0000101111 : logcos2 = mux_in_cos47;
        10'b0000110000 : logcos2 = mux_in_cos48;
        10'b0000110001 : logcos2 = mux_in_cos49;
        10'b0000110010 : logcos2 = mux_in_cos50;
        10'b0000110011 : logcos2 = mux_in_cos51;
        10'b0000110100 : logcos2 = mux_in_cos52;
        10'b0000110101 : logcos2 = mux_in_cos53;
        10'b0000110110 : logcos2 = mux_in_cos54;
        10'b0000110111 : logcos2 = mux_in_cos55;
        10'b0000111000 : logcos2 = mux_in_cos56;
        10'b0000111001 : logcos2 = mux_in_cos57;
        10'b0000111010 : logcos2 = mux_in_cos58;
        10'b0000111011 : logcos2 = mux_in_cos59;
        10'b0000111100 : logcos2 = mux_in_cos60;
        10'b0000111101 : logcos2 = mux_in_cos61;
        10'b0000111110 : logcos2 = mux_in_cos62;
        10'b0000111111 : logcos2 = mux_in_cos63;
        10'b0001000000 : logcos2 = mux_in_cos64;
        10'b0001000001 : logcos2 = mux_in_cos65;
        10'b0001000010 : logcos2 = mux_in_cos66;
        10'b0001000011 : logcos2 = mux_in_cos67;
        10'b0001000100 : logcos2 = mux_in_cos68;
        10'b0001000101 : logcos2 = mux_in_cos69;
        10'b0001000110 : logcos2 = mux_in_cos70;
        10'b0001000111 : logcos2 = mux_in_cos71;
        10'b0001001000 : logcos2 = mux_in_cos72;
        10'b0001001001 : logcos2 = mux_in_cos73;
        10'b0001001010 : logcos2 = mux_in_cos74;
        10'b0001001011 : logcos2 = mux_in_cos75;
        10'b0001001100 : logcos2 = mux_in_cos76;
        10'b0001001101 : logcos2 = mux_in_cos77;
        10'b0001001110 : logcos2 = mux_in_cos78;
        10'b0001001111 : logcos2 = mux_in_cos79;
        10'b0001010000 : logcos2 = mux_in_cos80;
        10'b0001010001 : logcos2 = mux_in_cos81;
        10'b0001010010 : logcos2 = mux_in_cos82;
        10'b0001010011 : logcos2 = mux_in_cos83;
        10'b0001010100 : logcos2 = mux_in_cos84;
        10'b0001010101 : logcos2 = mux_in_cos85;
        10'b0001010110 : logcos2 = mux_in_cos86;
        10'b0001010111 : logcos2 = mux_in_cos87;
        10'b0001011000 : logcos2 = mux_in_cos88;
        10'b0001011001 : logcos2 = mux_in_cos89;
        10'b0001011010 : logcos2 = mux_in_cos90;
        10'b0001011011 : logcos2 = mux_in_cos91;
        10'b0001011100 : logcos2 = mux_in_cos92;
        10'b0001011101 : logcos2 = mux_in_cos93;
        10'b0001011110 : logcos2 = mux_in_cos94;
        10'b0001011111 : logcos2 = mux_in_cos95;
        10'b0001100000 : logcos2 = mux_in_cos96;
        10'b0001100001 : logcos2 = mux_in_cos97;
        10'b0001100010 : logcos2 = mux_in_cos98;
        10'b0001100011 : logcos2 = mux_in_cos99;
        10'b0001100100 : logcos2 = mux_in_cos100;
        10'b0001100101 : logcos2 = mux_in_cos101;
        10'b0001100110 : logcos2 = mux_in_cos102;
        10'b0001100111 : logcos2 = mux_in_cos103;
        10'b0001101000 : logcos2 = mux_in_cos104;
        10'b0001101001 : logcos2 = mux_in_cos105;
        10'b0001101010 : logcos2 = mux_in_cos106;
        10'b0001101011 : logcos2 = mux_in_cos107;
        10'b0001101100 : logcos2 = mux_in_cos108;
        10'b0001101101 : logcos2 = mux_in_cos109;
        10'b0001101110 : logcos2 = mux_in_cos110;
        10'b0001101111 : logcos2 = mux_in_cos111;
        10'b0001110000 : logcos2 = mux_in_cos112;
        10'b0001110001 : logcos2 = mux_in_cos113;
        10'b0001110010 : logcos2 = mux_in_cos114;
        10'b0001110011 : logcos2 = mux_in_cos115;
        10'b0001110100 : logcos2 = mux_in_cos116;
        10'b0001110101 : logcos2 = mux_in_cos117;
        10'b0001110110 : logcos2 = mux_in_cos118;
        10'b0001110111 : logcos2 = mux_in_cos119;
        10'b0001111000 : logcos2 = mux_in_cos120;
        10'b0001111001 : logcos2 = mux_in_cos121;
        10'b0001111010 : logcos2 = mux_in_cos122;
        10'b0001111011 : logcos2 = mux_in_cos123;
        10'b0001111100 : logcos2 = mux_in_cos124;
        10'b0001111101 : logcos2 = mux_in_cos125;
        10'b0001111110 : logcos2 = mux_in_cos126;
        10'b0001111111 : logcos2 = mux_in_cos127;
        10'b0010000000 : logcos2 = mux_in_cos128;
        10'b0010000001 : logcos2 = mux_in_cos129;
        10'b0010000010 : logcos2 = mux_in_cos130;
        10'b0010000011 : logcos2 = mux_in_cos131;
        10'b0010000100 : logcos2 = mux_in_cos132;
        10'b0010000101 : logcos2 = mux_in_cos133;
        10'b0010000110 : logcos2 = mux_in_cos134;
        10'b0010000111 : logcos2 = mux_in_cos135;
        10'b0010001000 : logcos2 = mux_in_cos136;
        10'b0010001001 : logcos2 = mux_in_cos137;
        10'b0010001010 : logcos2 = mux_in_cos138;
        10'b0010001011 : logcos2 = mux_in_cos139;
        10'b0010001100 : logcos2 = mux_in_cos140;
        10'b0010001101 : logcos2 = mux_in_cos141;
        10'b0010001110 : logcos2 = mux_in_cos142;
        10'b0010001111 : logcos2 = mux_in_cos143;
        10'b0010010000 : logcos2 = mux_in_cos144;
        10'b0010010001 : logcos2 = mux_in_cos145;
        10'b0010010010 : logcos2 = mux_in_cos146;
        10'b0010010011 : logcos2 = mux_in_cos147;
        10'b0010010100 : logcos2 = mux_in_cos148;
        10'b0010010101 : logcos2 = mux_in_cos149;
        10'b0010010110 : logcos2 = mux_in_cos150;
        10'b0010010111 : logcos2 = mux_in_cos151;
        10'b0010011000 : logcos2 = mux_in_cos152;
        10'b0010011001 : logcos2 = mux_in_cos153;
        10'b0010011010 : logcos2 = mux_in_cos154;
        10'b0010011011 : logcos2 = mux_in_cos155;
        10'b0010011100 : logcos2 = mux_in_cos156;
        10'b0010011101 : logcos2 = mux_in_cos157;
        10'b0010011110 : logcos2 = mux_in_cos158;
        10'b0010011111 : logcos2 = mux_in_cos159;
        10'b0010100000 : logcos2 = mux_in_cos160;
        10'b0010100001 : logcos2 = mux_in_cos161;
        10'b0010100010 : logcos2 = mux_in_cos162;
        10'b0010100011 : logcos2 = mux_in_cos163;
        10'b0010100100 : logcos2 = mux_in_cos164;
        10'b0010100101 : logcos2 = mux_in_cos165;
        10'b0010100110 : logcos2 = mux_in_cos166;
        10'b0010100111 : logcos2 = mux_in_cos167;
        10'b0010101000 : logcos2 = mux_in_cos168;
        10'b0010101001 : logcos2 = mux_in_cos169;
        10'b0010101010 : logcos2 = mux_in_cos170;
        10'b0010101011 : logcos2 = mux_in_cos171;
        10'b0010101100 : logcos2 = mux_in_cos172;
        10'b0010101101 : logcos2 = mux_in_cos173;
        10'b0010101110 : logcos2 = mux_in_cos174;
        10'b0010101111 : logcos2 = mux_in_cos175;
        10'b0010110000 : logcos2 = mux_in_cos176;
        10'b0010110001 : logcos2 = mux_in_cos177;
        10'b0010110010 : logcos2 = mux_in_cos178;
        10'b0010110011 : logcos2 = mux_in_cos179;
        10'b0010110100 : logcos2 = mux_in_cos180;
        10'b0010110101 : logcos2 = mux_in_cos181;
        10'b0010110110 : logcos2 = mux_in_cos182;
        10'b0010110111 : logcos2 = mux_in_cos183;
        10'b0010111000 : logcos2 = mux_in_cos184;
        10'b0010111001 : logcos2 = mux_in_cos185;
        10'b0010111010 : logcos2 = mux_in_cos186;
        10'b0010111011 : logcos2 = mux_in_cos187;
        10'b0010111100 : logcos2 = mux_in_cos188;
        10'b0010111101 : logcos2 = mux_in_cos189;
        10'b0010111110 : logcos2 = mux_in_cos190;
        10'b0010111111 : logcos2 = mux_in_cos191;
        10'b0011000000 : logcos2 = mux_in_cos192;
        10'b0011000001 : logcos2 = mux_in_cos193;
        10'b0011000010 : logcos2 = mux_in_cos194;
        10'b0011000011 : logcos2 = mux_in_cos195;
        10'b0011000100 : logcos2 = mux_in_cos196;
        10'b0011000101 : logcos2 = mux_in_cos197;
        10'b0011000110 : logcos2 = mux_in_cos198;
        10'b0011000111 : logcos2 = mux_in_cos199;
        10'b0011001000 : logcos2 = mux_in_cos200;
        10'b0011001001 : logcos2 = mux_in_cos201;
        10'b0011001010 : logcos2 = mux_in_cos202;
        10'b0011001011 : logcos2 = mux_in_cos203;
        10'b0011001100 : logcos2 = mux_in_cos204;
        10'b0011001101 : logcos2 = mux_in_cos205;
        10'b0011001110 : logcos2 = mux_in_cos206;
        10'b0011001111 : logcos2 = mux_in_cos207;
        10'b0011010000 : logcos2 = mux_in_cos208;
        10'b0011010001 : logcos2 = mux_in_cos209;
        10'b0011010010 : logcos2 = mux_in_cos210;
        10'b0011010011 : logcos2 = mux_in_cos211;
        10'b0011010100 : logcos2 = mux_in_cos212;
        10'b0011010101 : logcos2 = mux_in_cos213;
        10'b0011010110 : logcos2 = mux_in_cos214;
        10'b0011010111 : logcos2 = mux_in_cos215;
        10'b0011011000 : logcos2 = mux_in_cos216;
        10'b0011011001 : logcos2 = mux_in_cos217;
        10'b0011011010 : logcos2 = mux_in_cos218;
        10'b0011011011 : logcos2 = mux_in_cos219;
        10'b0011011100 : logcos2 = mux_in_cos220;
        10'b0011011101 : logcos2 = mux_in_cos221;
        10'b0011011110 : logcos2 = mux_in_cos222;
        10'b0011011111 : logcos2 = mux_in_cos223;
        10'b0011100000 : logcos2 = mux_in_cos224;
        10'b0011100001 : logcos2 = mux_in_cos225;
        10'b0011100010 : logcos2 = mux_in_cos226;
        10'b0011100011 : logcos2 = mux_in_cos227;
        10'b0011100100 : logcos2 = mux_in_cos228;
        10'b0011100101 : logcos2 = mux_in_cos229;
        10'b0011100110 : logcos2 = mux_in_cos230;
        10'b0011100111 : logcos2 = mux_in_cos231;
        10'b0011101000 : logcos2 = mux_in_cos232;
        10'b0011101001 : logcos2 = mux_in_cos233;
        10'b0011101010 : logcos2 = mux_in_cos234;
        10'b0011101011 : logcos2 = mux_in_cos235;
        10'b0011101100 : logcos2 = mux_in_cos236;
        10'b0011101101 : logcos2 = mux_in_cos237;
        10'b0011101110 : logcos2 = mux_in_cos238;
        10'b0011101111 : logcos2 = mux_in_cos239;
        10'b0011110000 : logcos2 = mux_in_cos240;
        10'b0011110001 : logcos2 = mux_in_cos241;
        10'b0011110010 : logcos2 = mux_in_cos242;
        10'b0011110011 : logcos2 = mux_in_cos243;
        10'b0011110100 : logcos2 = mux_in_cos244;
        10'b0011110101 : logcos2 = mux_in_cos245;
        10'b0011110110 : logcos2 = mux_in_cos246;
        10'b0011110111 : logcos2 = mux_in_cos247;
        10'b0011111000 : logcos2 = mux_in_cos248;
        10'b0011111001 : logcos2 = mux_in_cos249;
        10'b0011111010 : logcos2 = mux_in_cos250;
        10'b0011111011 : logcos2 = mux_in_cos251;
        10'b0011111100 : logcos2 = mux_in_cos252;
        10'b0011111101 : logcos2 = mux_in_cos253;
        10'b0011111110 : logcos2 = mux_in_cos254;
        10'b0011111111 : logcos2 = mux_in_cos255;
        10'b0100000000 : logcos2 = mux_in_cos256;
        10'b0100000001 : logcos2 = mux_in_cos257;
        10'b0100000010 : logcos2 = mux_in_cos258;
        10'b0100000011 : logcos2 = mux_in_cos259;
        10'b0100000100 : logcos2 = mux_in_cos260;
        10'b0100000101 : logcos2 = mux_in_cos261;
        10'b0100000110 : logcos2 = mux_in_cos262;
        10'b0100000111 : logcos2 = mux_in_cos263;
        10'b0100001000 : logcos2 = mux_in_cos264;
        10'b0100001001 : logcos2 = mux_in_cos265;
        10'b0100001010 : logcos2 = mux_in_cos266;
        10'b0100001011 : logcos2 = mux_in_cos267;
        10'b0100001100 : logcos2 = mux_in_cos268;
        10'b0100001101 : logcos2 = mux_in_cos269;
        10'b0100001110 : logcos2 = mux_in_cos270;
        10'b0100001111 : logcos2 = mux_in_cos271;
        10'b0100010000 : logcos2 = mux_in_cos272;
        10'b0100010001 : logcos2 = mux_in_cos273;
        10'b0100010010 : logcos2 = mux_in_cos274;
        10'b0100010011 : logcos2 = mux_in_cos275;
        10'b0100010100 : logcos2 = mux_in_cos276;
        10'b0100010101 : logcos2 = mux_in_cos277;
        10'b0100010110 : logcos2 = mux_in_cos278;
        10'b0100010111 : logcos2 = mux_in_cos279;
        10'b0100011000 : logcos2 = mux_in_cos280;
        10'b0100011001 : logcos2 = mux_in_cos281;
        10'b0100011010 : logcos2 = mux_in_cos282;
        10'b0100011011 : logcos2 = mux_in_cos283;
        10'b0100011100 : logcos2 = mux_in_cos284;
        10'b0100011101 : logcos2 = mux_in_cos285;
        10'b0100011110 : logcos2 = mux_in_cos286;
        10'b0100011111 : logcos2 = mux_in_cos287;
        10'b0100100000 : logcos2 = mux_in_cos288;
        10'b0100100001 : logcos2 = mux_in_cos289;
        10'b0100100010 : logcos2 = mux_in_cos290;
        10'b0100100011 : logcos2 = mux_in_cos291;
        10'b0100100100 : logcos2 = mux_in_cos292;
        10'b0100100101 : logcos2 = mux_in_cos293;
        10'b0100100110 : logcos2 = mux_in_cos294;
        10'b0100100111 : logcos2 = mux_in_cos295;
        10'b0100101000 : logcos2 = mux_in_cos296;
        10'b0100101001 : logcos2 = mux_in_cos297;
        10'b0100101010 : logcos2 = mux_in_cos298;
        10'b0100101011 : logcos2 = mux_in_cos299;
        10'b0100101100 : logcos2 = mux_in_cos300;
        10'b0100101101 : logcos2 = mux_in_cos301;
        10'b0100101110 : logcos2 = mux_in_cos302;
        10'b0100101111 : logcos2 = mux_in_cos303;
        10'b0100110000 : logcos2 = mux_in_cos304;
        10'b0100110001 : logcos2 = mux_in_cos305;
        10'b0100110010 : logcos2 = mux_in_cos306;
        10'b0100110011 : logcos2 = mux_in_cos307;
        10'b0100110100 : logcos2 = mux_in_cos308;
        10'b0100110101 : logcos2 = mux_in_cos309;
        10'b0100110110 : logcos2 = mux_in_cos310;
        10'b0100110111 : logcos2 = mux_in_cos311;
        10'b0100111000 : logcos2 = mux_in_cos312;
        10'b0100111001 : logcos2 = mux_in_cos313;
        10'b0100111010 : logcos2 = mux_in_cos314;
        10'b0100111011 : logcos2 = mux_in_cos315;
        10'b0100111100 : logcos2 = mux_in_cos316;
        10'b0100111101 : logcos2 = mux_in_cos317;
        10'b0100111110 : logcos2 = mux_in_cos318;
        10'b0100111111 : logcos2 = mux_in_cos319;
        10'b0101000000 : logcos2 = mux_in_cos320;
        10'b0101000001 : logcos2 = mux_in_cos321;
        10'b0101000010 : logcos2 = mux_in_cos322;
        10'b0101000011 : logcos2 = mux_in_cos323;
        10'b0101000100 : logcos2 = mux_in_cos324;
        10'b0101000101 : logcos2 = mux_in_cos325;
        10'b0101000110 : logcos2 = mux_in_cos326;
        10'b0101000111 : logcos2 = mux_in_cos327;
        10'b0101001000 : logcos2 = mux_in_cos328;
        10'b0101001001 : logcos2 = mux_in_cos329;
        10'b0101001010 : logcos2 = mux_in_cos330;
        10'b0101001011 : logcos2 = mux_in_cos331;
        10'b0101001100 : logcos2 = mux_in_cos332;
        10'b0101001101 : logcos2 = mux_in_cos333;
        10'b0101001110 : logcos2 = mux_in_cos334;
        10'b0101001111 : logcos2 = mux_in_cos335;
        10'b0101010000 : logcos2 = mux_in_cos336;
        10'b0101010001 : logcos2 = mux_in_cos337;
        10'b0101010010 : logcos2 = mux_in_cos338;
        10'b0101010011 : logcos2 = mux_in_cos339;
        10'b0101010100 : logcos2 = mux_in_cos340;
        10'b0101010101 : logcos2 = mux_in_cos341;
        10'b0101010110 : logcos2 = mux_in_cos342;
        10'b0101010111 : logcos2 = mux_in_cos343;
        10'b0101011000 : logcos2 = mux_in_cos344;
        10'b0101011001 : logcos2 = mux_in_cos345;
        10'b0101011010 : logcos2 = mux_in_cos346;
        10'b0101011011 : logcos2 = mux_in_cos347;
        10'b0101011100 : logcos2 = mux_in_cos348;
        10'b0101011101 : logcos2 = mux_in_cos349;
        10'b0101011110 : logcos2 = mux_in_cos350;
        10'b0101011111 : logcos2 = mux_in_cos351;
        10'b0101100000 : logcos2 = mux_in_cos352;
        10'b0101100001 : logcos2 = mux_in_cos353;
        10'b0101100010 : logcos2 = mux_in_cos354;
        10'b0101100011 : logcos2 = mux_in_cos355;
        10'b0101100100 : logcos2 = mux_in_cos356;
        10'b0101100101 : logcos2 = mux_in_cos357;
        10'b0101100110 : logcos2 = mux_in_cos358;
        10'b0101100111 : logcos2 = mux_in_cos359;
        10'b0101101000 : logcos2 = mux_in_cos360;
        10'b0101101001 : logcos2 = mux_in_cos361;
        10'b0101101010 : logcos2 = mux_in_cos362;
        10'b0101101011 : logcos2 = mux_in_cos363;
        10'b0101101100 : logcos2 = mux_in_cos364;
        10'b0101101101 : logcos2 = mux_in_cos365;
        10'b0101101110 : logcos2 = mux_in_cos366;
        10'b0101101111 : logcos2 = mux_in_cos367;
        10'b0101110000 : logcos2 = mux_in_cos368;
        10'b0101110001 : logcos2 = mux_in_cos369;
        10'b0101110010 : logcos2 = mux_in_cos370;
        10'b0101110011 : logcos2 = mux_in_cos371;
        10'b0101110100 : logcos2 = mux_in_cos372;
        10'b0101110101 : logcos2 = mux_in_cos373;
        10'b0101110110 : logcos2 = mux_in_cos374;
        10'b0101110111 : logcos2 = mux_in_cos375;
        10'b0101111000 : logcos2 = mux_in_cos376;
        10'b0101111001 : logcos2 = mux_in_cos377;
        10'b0101111010 : logcos2 = mux_in_cos378;
        10'b0101111011 : logcos2 = mux_in_cos379;
        10'b0101111100 : logcos2 = mux_in_cos380;
        10'b0101111101 : logcos2 = mux_in_cos381;
        10'b0101111110 : logcos2 = mux_in_cos382;
        10'b0101111111 : logcos2 = mux_in_cos383;
        10'b0110000000 : logcos2 = mux_in_cos384;
        10'b0110000001 : logcos2 = mux_in_cos385;
        10'b0110000010 : logcos2 = mux_in_cos386;
        10'b0110000011 : logcos2 = mux_in_cos387;
        10'b0110000100 : logcos2 = mux_in_cos388;
        10'b0110000101 : logcos2 = mux_in_cos389;
        10'b0110000110 : logcos2 = mux_in_cos390;
        10'b0110000111 : logcos2 = mux_in_cos391;
        10'b0110001000 : logcos2 = mux_in_cos392;
        10'b0110001001 : logcos2 = mux_in_cos393;
        10'b0110001010 : logcos2 = mux_in_cos394;
        10'b0110001011 : logcos2 = mux_in_cos395;
        10'b0110001100 : logcos2 = mux_in_cos396;
        10'b0110001101 : logcos2 = mux_in_cos397;
        10'b0110001110 : logcos2 = mux_in_cos398;
        10'b0110001111 : logcos2 = mux_in_cos399;
        10'b0110010000 : logcos2 = mux_in_cos400;
        10'b0110010001 : logcos2 = mux_in_cos401;
        10'b0110010010 : logcos2 = mux_in_cos402;
        10'b0110010011 : logcos2 = mux_in_cos403;
        10'b0110010100 : logcos2 = mux_in_cos404;
        10'b0110010101 : logcos2 = mux_in_cos405;
        10'b0110010110 : logcos2 = mux_in_cos406;
        10'b0110010111 : logcos2 = mux_in_cos407;
        10'b0110011000 : logcos2 = mux_in_cos408;
        10'b0110011001 : logcos2 = mux_in_cos409;
        10'b0110011010 : logcos2 = mux_in_cos410;
        10'b0110011011 : logcos2 = mux_in_cos411;
        10'b0110011100 : logcos2 = mux_in_cos412;
        10'b0110011101 : logcos2 = mux_in_cos413;
        10'b0110011110 : logcos2 = mux_in_cos414;
        10'b0110011111 : logcos2 = mux_in_cos415;
        10'b0110100000 : logcos2 = mux_in_cos416;
        10'b0110100001 : logcos2 = mux_in_cos417;
        10'b0110100010 : logcos2 = mux_in_cos418;
        10'b0110100011 : logcos2 = mux_in_cos419;
        10'b0110100100 : logcos2 = mux_in_cos420;
        10'b0110100101 : logcos2 = mux_in_cos421;
        10'b0110100110 : logcos2 = mux_in_cos422;
        10'b0110100111 : logcos2 = mux_in_cos423;
        10'b0110101000 : logcos2 = mux_in_cos424;
        10'b0110101001 : logcos2 = mux_in_cos425;
        10'b0110101010 : logcos2 = mux_in_cos426;
        10'b0110101011 : logcos2 = mux_in_cos427;
        10'b0110101100 : logcos2 = mux_in_cos428;
        10'b0110101101 : logcos2 = mux_in_cos429;
        10'b0110101110 : logcos2 = mux_in_cos430;
        10'b0110101111 : logcos2 = mux_in_cos431;
        10'b0110110000 : logcos2 = mux_in_cos432;
        10'b0110110001 : logcos2 = mux_in_cos433;
        10'b0110110010 : logcos2 = mux_in_cos434;
        10'b0110110011 : logcos2 = mux_in_cos435;
        10'b0110110100 : logcos2 = mux_in_cos436;
        10'b0110110101 : logcos2 = mux_in_cos437;
        10'b0110110110 : logcos2 = mux_in_cos438;
        10'b0110110111 : logcos2 = mux_in_cos439;
        10'b0110111000 : logcos2 = mux_in_cos440;
        10'b0110111001 : logcos2 = mux_in_cos441;
        10'b0110111010 : logcos2 = mux_in_cos442;
        10'b0110111011 : logcos2 = mux_in_cos443;
        10'b0110111100 : logcos2 = mux_in_cos444;
        10'b0110111101 : logcos2 = mux_in_cos445;
        10'b0110111110 : logcos2 = mux_in_cos446;
        10'b0110111111 : logcos2 = mux_in_cos447;
        10'b0111000000 : logcos2 = mux_in_cos448;
        10'b0111000001 : logcos2 = mux_in_cos449;
        10'b0111000010 : logcos2 = mux_in_cos450;
        10'b0111000011 : logcos2 = mux_in_cos451;
        10'b0111000100 : logcos2 = mux_in_cos452;
        10'b0111000101 : logcos2 = mux_in_cos453;
        10'b0111000110 : logcos2 = mux_in_cos454;
        10'b0111000111 : logcos2 = mux_in_cos455;
        10'b0111001000 : logcos2 = mux_in_cos456;
        10'b0111001001 : logcos2 = mux_in_cos457;
        10'b0111001010 : logcos2 = mux_in_cos458;
        10'b0111001011 : logcos2 = mux_in_cos459;
        10'b0111001100 : logcos2 = mux_in_cos460;
        10'b0111001101 : logcos2 = mux_in_cos461;
        10'b0111001110 : logcos2 = mux_in_cos462;
        10'b0111001111 : logcos2 = mux_in_cos463;
        10'b0111010000 : logcos2 = mux_in_cos464;
        10'b0111010001 : logcos2 = mux_in_cos465;
        10'b0111010010 : logcos2 = mux_in_cos466;
        10'b0111010011 : logcos2 = mux_in_cos467;
        10'b0111010100 : logcos2 = mux_in_cos468;
        10'b0111010101 : logcos2 = mux_in_cos469;
        10'b0111010110 : logcos2 = mux_in_cos470;
        10'b0111010111 : logcos2 = mux_in_cos471;
        10'b0111011000 : logcos2 = mux_in_cos472;
        10'b0111011001 : logcos2 = mux_in_cos473;
        10'b0111011010 : logcos2 = mux_in_cos474;
        10'b0111011011 : logcos2 = mux_in_cos475;
        10'b0111011100 : logcos2 = mux_in_cos476;
        10'b0111011101 : logcos2 = mux_in_cos477;
        10'b0111011110 : logcos2 = mux_in_cos478;
        10'b0111011111 : logcos2 = mux_in_cos479;
        10'b0111100000 : logcos2 = mux_in_cos480;
        10'b0111100001 : logcos2 = mux_in_cos481;
        10'b0111100010 : logcos2 = mux_in_cos482;
        10'b0111100011 : logcos2 = mux_in_cos483;
        10'b0111100100 : logcos2 = mux_in_cos484;
        10'b0111100101 : logcos2 = mux_in_cos485;
        10'b0111100110 : logcos2 = mux_in_cos486;
        10'b0111100111 : logcos2 = mux_in_cos487;
        10'b0111101000 : logcos2 = mux_in_cos488;
        10'b0111101001 : logcos2 = mux_in_cos489;
        10'b0111101010 : logcos2 = mux_in_cos490;
        10'b0111101011 : logcos2 = mux_in_cos491;
        10'b0111101100 : logcos2 = mux_in_cos492;
        10'b0111101101 : logcos2 = mux_in_cos493;
        10'b0111101110 : logcos2 = mux_in_cos494;
        10'b0111101111 : logcos2 = mux_in_cos495;
        10'b0111110000 : logcos2 = mux_in_cos496;
        10'b0111110001 : logcos2 = mux_in_cos497;
        10'b0111110010 : logcos2 = mux_in_cos498;
        10'b0111110011 : logcos2 = mux_in_cos499;
        10'b0111110100 : logcos2 = mux_in_cos500;
        10'b0111110101 : logcos2 = mux_in_cos501;
        10'b0111110110 : logcos2 = mux_in_cos502;
        10'b0111110111 : logcos2 = mux_in_cos503;
        10'b0111111000 : logcos2 = mux_in_cos504;
        10'b0111111001 : logcos2 = mux_in_cos505;
        10'b0111111010 : logcos2 = mux_in_cos506;
        10'b0111111011 : logcos2 = mux_in_cos507;
        10'b0111111100 : logcos2 = mux_in_cos508;
        10'b0111111101 : logcos2 = mux_in_cos509;
        10'b0111111110 : logcos2 = mux_in_cos510;
        10'b0111111111 : logcos2 = mux_in_cos511;
        10'b1000000000 : logcos2 = mux_in_cos512;
        default: logcos2 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in3)
        10'b0000000000 : logcos3 = mux_in_cos0;
        10'b0000000001 : logcos3 = mux_in_cos1;
        10'b0000000010 : logcos3 = mux_in_cos2;
        10'b0000000011 : logcos3 = mux_in_cos3;
        10'b0000000100 : logcos3 = mux_in_cos4;
        10'b0000000101 : logcos3 = mux_in_cos5;
        10'b0000000110 : logcos3 = mux_in_cos6;
        10'b0000000111 : logcos3 = mux_in_cos7;
        10'b0000001000 : logcos3 = mux_in_cos8;
        10'b0000001001 : logcos3 = mux_in_cos9;
        10'b0000001010 : logcos3 = mux_in_cos10;
        10'b0000001011 : logcos3 = mux_in_cos11;
        10'b0000001100 : logcos3 = mux_in_cos12;
        10'b0000001101 : logcos3 = mux_in_cos13;
        10'b0000001110 : logcos3 = mux_in_cos14;
        10'b0000001111 : logcos3 = mux_in_cos15;
        10'b0000010000 : logcos3 = mux_in_cos16;
        10'b0000010001 : logcos3 = mux_in_cos17;
        10'b0000010010 : logcos3 = mux_in_cos18;
        10'b0000010011 : logcos3 = mux_in_cos19;
        10'b0000010100 : logcos3 = mux_in_cos20;
        10'b0000010101 : logcos3 = mux_in_cos21;
        10'b0000010110 : logcos3 = mux_in_cos22;
        10'b0000010111 : logcos3 = mux_in_cos23;
        10'b0000011000 : logcos3 = mux_in_cos24;
        10'b0000011001 : logcos3 = mux_in_cos25;
        10'b0000011010 : logcos3 = mux_in_cos26;
        10'b0000011011 : logcos3 = mux_in_cos27;
        10'b0000011100 : logcos3 = mux_in_cos28;
        10'b0000011101 : logcos3 = mux_in_cos29;
        10'b0000011110 : logcos3 = mux_in_cos30;
        10'b0000011111 : logcos3 = mux_in_cos31;
        10'b0000100000 : logcos3 = mux_in_cos32;
        10'b0000100001 : logcos3 = mux_in_cos33;
        10'b0000100010 : logcos3 = mux_in_cos34;
        10'b0000100011 : logcos3 = mux_in_cos35;
        10'b0000100100 : logcos3 = mux_in_cos36;
        10'b0000100101 : logcos3 = mux_in_cos37;
        10'b0000100110 : logcos3 = mux_in_cos38;
        10'b0000100111 : logcos3 = mux_in_cos39;
        10'b0000101000 : logcos3 = mux_in_cos40;
        10'b0000101001 : logcos3 = mux_in_cos41;
        10'b0000101010 : logcos3 = mux_in_cos42;
        10'b0000101011 : logcos3 = mux_in_cos43;
        10'b0000101100 : logcos3 = mux_in_cos44;
        10'b0000101101 : logcos3 = mux_in_cos45;
        10'b0000101110 : logcos3 = mux_in_cos46;
        10'b0000101111 : logcos3 = mux_in_cos47;
        10'b0000110000 : logcos3 = mux_in_cos48;
        10'b0000110001 : logcos3 = mux_in_cos49;
        10'b0000110010 : logcos3 = mux_in_cos50;
        10'b0000110011 : logcos3 = mux_in_cos51;
        10'b0000110100 : logcos3 = mux_in_cos52;
        10'b0000110101 : logcos3 = mux_in_cos53;
        10'b0000110110 : logcos3 = mux_in_cos54;
        10'b0000110111 : logcos3 = mux_in_cos55;
        10'b0000111000 : logcos3 = mux_in_cos56;
        10'b0000111001 : logcos3 = mux_in_cos57;
        10'b0000111010 : logcos3 = mux_in_cos58;
        10'b0000111011 : logcos3 = mux_in_cos59;
        10'b0000111100 : logcos3 = mux_in_cos60;
        10'b0000111101 : logcos3 = mux_in_cos61;
        10'b0000111110 : logcos3 = mux_in_cos62;
        10'b0000111111 : logcos3 = mux_in_cos63;
        10'b0001000000 : logcos3 = mux_in_cos64;
        10'b0001000001 : logcos3 = mux_in_cos65;
        10'b0001000010 : logcos3 = mux_in_cos66;
        10'b0001000011 : logcos3 = mux_in_cos67;
        10'b0001000100 : logcos3 = mux_in_cos68;
        10'b0001000101 : logcos3 = mux_in_cos69;
        10'b0001000110 : logcos3 = mux_in_cos70;
        10'b0001000111 : logcos3 = mux_in_cos71;
        10'b0001001000 : logcos3 = mux_in_cos72;
        10'b0001001001 : logcos3 = mux_in_cos73;
        10'b0001001010 : logcos3 = mux_in_cos74;
        10'b0001001011 : logcos3 = mux_in_cos75;
        10'b0001001100 : logcos3 = mux_in_cos76;
        10'b0001001101 : logcos3 = mux_in_cos77;
        10'b0001001110 : logcos3 = mux_in_cos78;
        10'b0001001111 : logcos3 = mux_in_cos79;
        10'b0001010000 : logcos3 = mux_in_cos80;
        10'b0001010001 : logcos3 = mux_in_cos81;
        10'b0001010010 : logcos3 = mux_in_cos82;
        10'b0001010011 : logcos3 = mux_in_cos83;
        10'b0001010100 : logcos3 = mux_in_cos84;
        10'b0001010101 : logcos3 = mux_in_cos85;
        10'b0001010110 : logcos3 = mux_in_cos86;
        10'b0001010111 : logcos3 = mux_in_cos87;
        10'b0001011000 : logcos3 = mux_in_cos88;
        10'b0001011001 : logcos3 = mux_in_cos89;
        10'b0001011010 : logcos3 = mux_in_cos90;
        10'b0001011011 : logcos3 = mux_in_cos91;
        10'b0001011100 : logcos3 = mux_in_cos92;
        10'b0001011101 : logcos3 = mux_in_cos93;
        10'b0001011110 : logcos3 = mux_in_cos94;
        10'b0001011111 : logcos3 = mux_in_cos95;
        10'b0001100000 : logcos3 = mux_in_cos96;
        10'b0001100001 : logcos3 = mux_in_cos97;
        10'b0001100010 : logcos3 = mux_in_cos98;
        10'b0001100011 : logcos3 = mux_in_cos99;
        10'b0001100100 : logcos3 = mux_in_cos100;
        10'b0001100101 : logcos3 = mux_in_cos101;
        10'b0001100110 : logcos3 = mux_in_cos102;
        10'b0001100111 : logcos3 = mux_in_cos103;
        10'b0001101000 : logcos3 = mux_in_cos104;
        10'b0001101001 : logcos3 = mux_in_cos105;
        10'b0001101010 : logcos3 = mux_in_cos106;
        10'b0001101011 : logcos3 = mux_in_cos107;
        10'b0001101100 : logcos3 = mux_in_cos108;
        10'b0001101101 : logcos3 = mux_in_cos109;
        10'b0001101110 : logcos3 = mux_in_cos110;
        10'b0001101111 : logcos3 = mux_in_cos111;
        10'b0001110000 : logcos3 = mux_in_cos112;
        10'b0001110001 : logcos3 = mux_in_cos113;
        10'b0001110010 : logcos3 = mux_in_cos114;
        10'b0001110011 : logcos3 = mux_in_cos115;
        10'b0001110100 : logcos3 = mux_in_cos116;
        10'b0001110101 : logcos3 = mux_in_cos117;
        10'b0001110110 : logcos3 = mux_in_cos118;
        10'b0001110111 : logcos3 = mux_in_cos119;
        10'b0001111000 : logcos3 = mux_in_cos120;
        10'b0001111001 : logcos3 = mux_in_cos121;
        10'b0001111010 : logcos3 = mux_in_cos122;
        10'b0001111011 : logcos3 = mux_in_cos123;
        10'b0001111100 : logcos3 = mux_in_cos124;
        10'b0001111101 : logcos3 = mux_in_cos125;
        10'b0001111110 : logcos3 = mux_in_cos126;
        10'b0001111111 : logcos3 = mux_in_cos127;
        10'b0010000000 : logcos3 = mux_in_cos128;
        10'b0010000001 : logcos3 = mux_in_cos129;
        10'b0010000010 : logcos3 = mux_in_cos130;
        10'b0010000011 : logcos3 = mux_in_cos131;
        10'b0010000100 : logcos3 = mux_in_cos132;
        10'b0010000101 : logcos3 = mux_in_cos133;
        10'b0010000110 : logcos3 = mux_in_cos134;
        10'b0010000111 : logcos3 = mux_in_cos135;
        10'b0010001000 : logcos3 = mux_in_cos136;
        10'b0010001001 : logcos3 = mux_in_cos137;
        10'b0010001010 : logcos3 = mux_in_cos138;
        10'b0010001011 : logcos3 = mux_in_cos139;
        10'b0010001100 : logcos3 = mux_in_cos140;
        10'b0010001101 : logcos3 = mux_in_cos141;
        10'b0010001110 : logcos3 = mux_in_cos142;
        10'b0010001111 : logcos3 = mux_in_cos143;
        10'b0010010000 : logcos3 = mux_in_cos144;
        10'b0010010001 : logcos3 = mux_in_cos145;
        10'b0010010010 : logcos3 = mux_in_cos146;
        10'b0010010011 : logcos3 = mux_in_cos147;
        10'b0010010100 : logcos3 = mux_in_cos148;
        10'b0010010101 : logcos3 = mux_in_cos149;
        10'b0010010110 : logcos3 = mux_in_cos150;
        10'b0010010111 : logcos3 = mux_in_cos151;
        10'b0010011000 : logcos3 = mux_in_cos152;
        10'b0010011001 : logcos3 = mux_in_cos153;
        10'b0010011010 : logcos3 = mux_in_cos154;
        10'b0010011011 : logcos3 = mux_in_cos155;
        10'b0010011100 : logcos3 = mux_in_cos156;
        10'b0010011101 : logcos3 = mux_in_cos157;
        10'b0010011110 : logcos3 = mux_in_cos158;
        10'b0010011111 : logcos3 = mux_in_cos159;
        10'b0010100000 : logcos3 = mux_in_cos160;
        10'b0010100001 : logcos3 = mux_in_cos161;
        10'b0010100010 : logcos3 = mux_in_cos162;
        10'b0010100011 : logcos3 = mux_in_cos163;
        10'b0010100100 : logcos3 = mux_in_cos164;
        10'b0010100101 : logcos3 = mux_in_cos165;
        10'b0010100110 : logcos3 = mux_in_cos166;
        10'b0010100111 : logcos3 = mux_in_cos167;
        10'b0010101000 : logcos3 = mux_in_cos168;
        10'b0010101001 : logcos3 = mux_in_cos169;
        10'b0010101010 : logcos3 = mux_in_cos170;
        10'b0010101011 : logcos3 = mux_in_cos171;
        10'b0010101100 : logcos3 = mux_in_cos172;
        10'b0010101101 : logcos3 = mux_in_cos173;
        10'b0010101110 : logcos3 = mux_in_cos174;
        10'b0010101111 : logcos3 = mux_in_cos175;
        10'b0010110000 : logcos3 = mux_in_cos176;
        10'b0010110001 : logcos3 = mux_in_cos177;
        10'b0010110010 : logcos3 = mux_in_cos178;
        10'b0010110011 : logcos3 = mux_in_cos179;
        10'b0010110100 : logcos3 = mux_in_cos180;
        10'b0010110101 : logcos3 = mux_in_cos181;
        10'b0010110110 : logcos3 = mux_in_cos182;
        10'b0010110111 : logcos3 = mux_in_cos183;
        10'b0010111000 : logcos3 = mux_in_cos184;
        10'b0010111001 : logcos3 = mux_in_cos185;
        10'b0010111010 : logcos3 = mux_in_cos186;
        10'b0010111011 : logcos3 = mux_in_cos187;
        10'b0010111100 : logcos3 = mux_in_cos188;
        10'b0010111101 : logcos3 = mux_in_cos189;
        10'b0010111110 : logcos3 = mux_in_cos190;
        10'b0010111111 : logcos3 = mux_in_cos191;
        10'b0011000000 : logcos3 = mux_in_cos192;
        10'b0011000001 : logcos3 = mux_in_cos193;
        10'b0011000010 : logcos3 = mux_in_cos194;
        10'b0011000011 : logcos3 = mux_in_cos195;
        10'b0011000100 : logcos3 = mux_in_cos196;
        10'b0011000101 : logcos3 = mux_in_cos197;
        10'b0011000110 : logcos3 = mux_in_cos198;
        10'b0011000111 : logcos3 = mux_in_cos199;
        10'b0011001000 : logcos3 = mux_in_cos200;
        10'b0011001001 : logcos3 = mux_in_cos201;
        10'b0011001010 : logcos3 = mux_in_cos202;
        10'b0011001011 : logcos3 = mux_in_cos203;
        10'b0011001100 : logcos3 = mux_in_cos204;
        10'b0011001101 : logcos3 = mux_in_cos205;
        10'b0011001110 : logcos3 = mux_in_cos206;
        10'b0011001111 : logcos3 = mux_in_cos207;
        10'b0011010000 : logcos3 = mux_in_cos208;
        10'b0011010001 : logcos3 = mux_in_cos209;
        10'b0011010010 : logcos3 = mux_in_cos210;
        10'b0011010011 : logcos3 = mux_in_cos211;
        10'b0011010100 : logcos3 = mux_in_cos212;
        10'b0011010101 : logcos3 = mux_in_cos213;
        10'b0011010110 : logcos3 = mux_in_cos214;
        10'b0011010111 : logcos3 = mux_in_cos215;
        10'b0011011000 : logcos3 = mux_in_cos216;
        10'b0011011001 : logcos3 = mux_in_cos217;
        10'b0011011010 : logcos3 = mux_in_cos218;
        10'b0011011011 : logcos3 = mux_in_cos219;
        10'b0011011100 : logcos3 = mux_in_cos220;
        10'b0011011101 : logcos3 = mux_in_cos221;
        10'b0011011110 : logcos3 = mux_in_cos222;
        10'b0011011111 : logcos3 = mux_in_cos223;
        10'b0011100000 : logcos3 = mux_in_cos224;
        10'b0011100001 : logcos3 = mux_in_cos225;
        10'b0011100010 : logcos3 = mux_in_cos226;
        10'b0011100011 : logcos3 = mux_in_cos227;
        10'b0011100100 : logcos3 = mux_in_cos228;
        10'b0011100101 : logcos3 = mux_in_cos229;
        10'b0011100110 : logcos3 = mux_in_cos230;
        10'b0011100111 : logcos3 = mux_in_cos231;
        10'b0011101000 : logcos3 = mux_in_cos232;
        10'b0011101001 : logcos3 = mux_in_cos233;
        10'b0011101010 : logcos3 = mux_in_cos234;
        10'b0011101011 : logcos3 = mux_in_cos235;
        10'b0011101100 : logcos3 = mux_in_cos236;
        10'b0011101101 : logcos3 = mux_in_cos237;
        10'b0011101110 : logcos3 = mux_in_cos238;
        10'b0011101111 : logcos3 = mux_in_cos239;
        10'b0011110000 : logcos3 = mux_in_cos240;
        10'b0011110001 : logcos3 = mux_in_cos241;
        10'b0011110010 : logcos3 = mux_in_cos242;
        10'b0011110011 : logcos3 = mux_in_cos243;
        10'b0011110100 : logcos3 = mux_in_cos244;
        10'b0011110101 : logcos3 = mux_in_cos245;
        10'b0011110110 : logcos3 = mux_in_cos246;
        10'b0011110111 : logcos3 = mux_in_cos247;
        10'b0011111000 : logcos3 = mux_in_cos248;
        10'b0011111001 : logcos3 = mux_in_cos249;
        10'b0011111010 : logcos3 = mux_in_cos250;
        10'b0011111011 : logcos3 = mux_in_cos251;
        10'b0011111100 : logcos3 = mux_in_cos252;
        10'b0011111101 : logcos3 = mux_in_cos253;
        10'b0011111110 : logcos3 = mux_in_cos254;
        10'b0011111111 : logcos3 = mux_in_cos255;
        10'b0100000000 : logcos3 = mux_in_cos256;
        10'b0100000001 : logcos3 = mux_in_cos257;
        10'b0100000010 : logcos3 = mux_in_cos258;
        10'b0100000011 : logcos3 = mux_in_cos259;
        10'b0100000100 : logcos3 = mux_in_cos260;
        10'b0100000101 : logcos3 = mux_in_cos261;
        10'b0100000110 : logcos3 = mux_in_cos262;
        10'b0100000111 : logcos3 = mux_in_cos263;
        10'b0100001000 : logcos3 = mux_in_cos264;
        10'b0100001001 : logcos3 = mux_in_cos265;
        10'b0100001010 : logcos3 = mux_in_cos266;
        10'b0100001011 : logcos3 = mux_in_cos267;
        10'b0100001100 : logcos3 = mux_in_cos268;
        10'b0100001101 : logcos3 = mux_in_cos269;
        10'b0100001110 : logcos3 = mux_in_cos270;
        10'b0100001111 : logcos3 = mux_in_cos271;
        10'b0100010000 : logcos3 = mux_in_cos272;
        10'b0100010001 : logcos3 = mux_in_cos273;
        10'b0100010010 : logcos3 = mux_in_cos274;
        10'b0100010011 : logcos3 = mux_in_cos275;
        10'b0100010100 : logcos3 = mux_in_cos276;
        10'b0100010101 : logcos3 = mux_in_cos277;
        10'b0100010110 : logcos3 = mux_in_cos278;
        10'b0100010111 : logcos3 = mux_in_cos279;
        10'b0100011000 : logcos3 = mux_in_cos280;
        10'b0100011001 : logcos3 = mux_in_cos281;
        10'b0100011010 : logcos3 = mux_in_cos282;
        10'b0100011011 : logcos3 = mux_in_cos283;
        10'b0100011100 : logcos3 = mux_in_cos284;
        10'b0100011101 : logcos3 = mux_in_cos285;
        10'b0100011110 : logcos3 = mux_in_cos286;
        10'b0100011111 : logcos3 = mux_in_cos287;
        10'b0100100000 : logcos3 = mux_in_cos288;
        10'b0100100001 : logcos3 = mux_in_cos289;
        10'b0100100010 : logcos3 = mux_in_cos290;
        10'b0100100011 : logcos3 = mux_in_cos291;
        10'b0100100100 : logcos3 = mux_in_cos292;
        10'b0100100101 : logcos3 = mux_in_cos293;
        10'b0100100110 : logcos3 = mux_in_cos294;
        10'b0100100111 : logcos3 = mux_in_cos295;
        10'b0100101000 : logcos3 = mux_in_cos296;
        10'b0100101001 : logcos3 = mux_in_cos297;
        10'b0100101010 : logcos3 = mux_in_cos298;
        10'b0100101011 : logcos3 = mux_in_cos299;
        10'b0100101100 : logcos3 = mux_in_cos300;
        10'b0100101101 : logcos3 = mux_in_cos301;
        10'b0100101110 : logcos3 = mux_in_cos302;
        10'b0100101111 : logcos3 = mux_in_cos303;
        10'b0100110000 : logcos3 = mux_in_cos304;
        10'b0100110001 : logcos3 = mux_in_cos305;
        10'b0100110010 : logcos3 = mux_in_cos306;
        10'b0100110011 : logcos3 = mux_in_cos307;
        10'b0100110100 : logcos3 = mux_in_cos308;
        10'b0100110101 : logcos3 = mux_in_cos309;
        10'b0100110110 : logcos3 = mux_in_cos310;
        10'b0100110111 : logcos3 = mux_in_cos311;
        10'b0100111000 : logcos3 = mux_in_cos312;
        10'b0100111001 : logcos3 = mux_in_cos313;
        10'b0100111010 : logcos3 = mux_in_cos314;
        10'b0100111011 : logcos3 = mux_in_cos315;
        10'b0100111100 : logcos3 = mux_in_cos316;
        10'b0100111101 : logcos3 = mux_in_cos317;
        10'b0100111110 : logcos3 = mux_in_cos318;
        10'b0100111111 : logcos3 = mux_in_cos319;
        10'b0101000000 : logcos3 = mux_in_cos320;
        10'b0101000001 : logcos3 = mux_in_cos321;
        10'b0101000010 : logcos3 = mux_in_cos322;
        10'b0101000011 : logcos3 = mux_in_cos323;
        10'b0101000100 : logcos3 = mux_in_cos324;
        10'b0101000101 : logcos3 = mux_in_cos325;
        10'b0101000110 : logcos3 = mux_in_cos326;
        10'b0101000111 : logcos3 = mux_in_cos327;
        10'b0101001000 : logcos3 = mux_in_cos328;
        10'b0101001001 : logcos3 = mux_in_cos329;
        10'b0101001010 : logcos3 = mux_in_cos330;
        10'b0101001011 : logcos3 = mux_in_cos331;
        10'b0101001100 : logcos3 = mux_in_cos332;
        10'b0101001101 : logcos3 = mux_in_cos333;
        10'b0101001110 : logcos3 = mux_in_cos334;
        10'b0101001111 : logcos3 = mux_in_cos335;
        10'b0101010000 : logcos3 = mux_in_cos336;
        10'b0101010001 : logcos3 = mux_in_cos337;
        10'b0101010010 : logcos3 = mux_in_cos338;
        10'b0101010011 : logcos3 = mux_in_cos339;
        10'b0101010100 : logcos3 = mux_in_cos340;
        10'b0101010101 : logcos3 = mux_in_cos341;
        10'b0101010110 : logcos3 = mux_in_cos342;
        10'b0101010111 : logcos3 = mux_in_cos343;
        10'b0101011000 : logcos3 = mux_in_cos344;
        10'b0101011001 : logcos3 = mux_in_cos345;
        10'b0101011010 : logcos3 = mux_in_cos346;
        10'b0101011011 : logcos3 = mux_in_cos347;
        10'b0101011100 : logcos3 = mux_in_cos348;
        10'b0101011101 : logcos3 = mux_in_cos349;
        10'b0101011110 : logcos3 = mux_in_cos350;
        10'b0101011111 : logcos3 = mux_in_cos351;
        10'b0101100000 : logcos3 = mux_in_cos352;
        10'b0101100001 : logcos3 = mux_in_cos353;
        10'b0101100010 : logcos3 = mux_in_cos354;
        10'b0101100011 : logcos3 = mux_in_cos355;
        10'b0101100100 : logcos3 = mux_in_cos356;
        10'b0101100101 : logcos3 = mux_in_cos357;
        10'b0101100110 : logcos3 = mux_in_cos358;
        10'b0101100111 : logcos3 = mux_in_cos359;
        10'b0101101000 : logcos3 = mux_in_cos360;
        10'b0101101001 : logcos3 = mux_in_cos361;
        10'b0101101010 : logcos3 = mux_in_cos362;
        10'b0101101011 : logcos3 = mux_in_cos363;
        10'b0101101100 : logcos3 = mux_in_cos364;
        10'b0101101101 : logcos3 = mux_in_cos365;
        10'b0101101110 : logcos3 = mux_in_cos366;
        10'b0101101111 : logcos3 = mux_in_cos367;
        10'b0101110000 : logcos3 = mux_in_cos368;
        10'b0101110001 : logcos3 = mux_in_cos369;
        10'b0101110010 : logcos3 = mux_in_cos370;
        10'b0101110011 : logcos3 = mux_in_cos371;
        10'b0101110100 : logcos3 = mux_in_cos372;
        10'b0101110101 : logcos3 = mux_in_cos373;
        10'b0101110110 : logcos3 = mux_in_cos374;
        10'b0101110111 : logcos3 = mux_in_cos375;
        10'b0101111000 : logcos3 = mux_in_cos376;
        10'b0101111001 : logcos3 = mux_in_cos377;
        10'b0101111010 : logcos3 = mux_in_cos378;
        10'b0101111011 : logcos3 = mux_in_cos379;
        10'b0101111100 : logcos3 = mux_in_cos380;
        10'b0101111101 : logcos3 = mux_in_cos381;
        10'b0101111110 : logcos3 = mux_in_cos382;
        10'b0101111111 : logcos3 = mux_in_cos383;
        10'b0110000000 : logcos3 = mux_in_cos384;
        10'b0110000001 : logcos3 = mux_in_cos385;
        10'b0110000010 : logcos3 = mux_in_cos386;
        10'b0110000011 : logcos3 = mux_in_cos387;
        10'b0110000100 : logcos3 = mux_in_cos388;
        10'b0110000101 : logcos3 = mux_in_cos389;
        10'b0110000110 : logcos3 = mux_in_cos390;
        10'b0110000111 : logcos3 = mux_in_cos391;
        10'b0110001000 : logcos3 = mux_in_cos392;
        10'b0110001001 : logcos3 = mux_in_cos393;
        10'b0110001010 : logcos3 = mux_in_cos394;
        10'b0110001011 : logcos3 = mux_in_cos395;
        10'b0110001100 : logcos3 = mux_in_cos396;
        10'b0110001101 : logcos3 = mux_in_cos397;
        10'b0110001110 : logcos3 = mux_in_cos398;
        10'b0110001111 : logcos3 = mux_in_cos399;
        10'b0110010000 : logcos3 = mux_in_cos400;
        10'b0110010001 : logcos3 = mux_in_cos401;
        10'b0110010010 : logcos3 = mux_in_cos402;
        10'b0110010011 : logcos3 = mux_in_cos403;
        10'b0110010100 : logcos3 = mux_in_cos404;
        10'b0110010101 : logcos3 = mux_in_cos405;
        10'b0110010110 : logcos3 = mux_in_cos406;
        10'b0110010111 : logcos3 = mux_in_cos407;
        10'b0110011000 : logcos3 = mux_in_cos408;
        10'b0110011001 : logcos3 = mux_in_cos409;
        10'b0110011010 : logcos3 = mux_in_cos410;
        10'b0110011011 : logcos3 = mux_in_cos411;
        10'b0110011100 : logcos3 = mux_in_cos412;
        10'b0110011101 : logcos3 = mux_in_cos413;
        10'b0110011110 : logcos3 = mux_in_cos414;
        10'b0110011111 : logcos3 = mux_in_cos415;
        10'b0110100000 : logcos3 = mux_in_cos416;
        10'b0110100001 : logcos3 = mux_in_cos417;
        10'b0110100010 : logcos3 = mux_in_cos418;
        10'b0110100011 : logcos3 = mux_in_cos419;
        10'b0110100100 : logcos3 = mux_in_cos420;
        10'b0110100101 : logcos3 = mux_in_cos421;
        10'b0110100110 : logcos3 = mux_in_cos422;
        10'b0110100111 : logcos3 = mux_in_cos423;
        10'b0110101000 : logcos3 = mux_in_cos424;
        10'b0110101001 : logcos3 = mux_in_cos425;
        10'b0110101010 : logcos3 = mux_in_cos426;
        10'b0110101011 : logcos3 = mux_in_cos427;
        10'b0110101100 : logcos3 = mux_in_cos428;
        10'b0110101101 : logcos3 = mux_in_cos429;
        10'b0110101110 : logcos3 = mux_in_cos430;
        10'b0110101111 : logcos3 = mux_in_cos431;
        10'b0110110000 : logcos3 = mux_in_cos432;
        10'b0110110001 : logcos3 = mux_in_cos433;
        10'b0110110010 : logcos3 = mux_in_cos434;
        10'b0110110011 : logcos3 = mux_in_cos435;
        10'b0110110100 : logcos3 = mux_in_cos436;
        10'b0110110101 : logcos3 = mux_in_cos437;
        10'b0110110110 : logcos3 = mux_in_cos438;
        10'b0110110111 : logcos3 = mux_in_cos439;
        10'b0110111000 : logcos3 = mux_in_cos440;
        10'b0110111001 : logcos3 = mux_in_cos441;
        10'b0110111010 : logcos3 = mux_in_cos442;
        10'b0110111011 : logcos3 = mux_in_cos443;
        10'b0110111100 : logcos3 = mux_in_cos444;
        10'b0110111101 : logcos3 = mux_in_cos445;
        10'b0110111110 : logcos3 = mux_in_cos446;
        10'b0110111111 : logcos3 = mux_in_cos447;
        10'b0111000000 : logcos3 = mux_in_cos448;
        10'b0111000001 : logcos3 = mux_in_cos449;
        10'b0111000010 : logcos3 = mux_in_cos450;
        10'b0111000011 : logcos3 = mux_in_cos451;
        10'b0111000100 : logcos3 = mux_in_cos452;
        10'b0111000101 : logcos3 = mux_in_cos453;
        10'b0111000110 : logcos3 = mux_in_cos454;
        10'b0111000111 : logcos3 = mux_in_cos455;
        10'b0111001000 : logcos3 = mux_in_cos456;
        10'b0111001001 : logcos3 = mux_in_cos457;
        10'b0111001010 : logcos3 = mux_in_cos458;
        10'b0111001011 : logcos3 = mux_in_cos459;
        10'b0111001100 : logcos3 = mux_in_cos460;
        10'b0111001101 : logcos3 = mux_in_cos461;
        10'b0111001110 : logcos3 = mux_in_cos462;
        10'b0111001111 : logcos3 = mux_in_cos463;
        10'b0111010000 : logcos3 = mux_in_cos464;
        10'b0111010001 : logcos3 = mux_in_cos465;
        10'b0111010010 : logcos3 = mux_in_cos466;
        10'b0111010011 : logcos3 = mux_in_cos467;
        10'b0111010100 : logcos3 = mux_in_cos468;
        10'b0111010101 : logcos3 = mux_in_cos469;
        10'b0111010110 : logcos3 = mux_in_cos470;
        10'b0111010111 : logcos3 = mux_in_cos471;
        10'b0111011000 : logcos3 = mux_in_cos472;
        10'b0111011001 : logcos3 = mux_in_cos473;
        10'b0111011010 : logcos3 = mux_in_cos474;
        10'b0111011011 : logcos3 = mux_in_cos475;
        10'b0111011100 : logcos3 = mux_in_cos476;
        10'b0111011101 : logcos3 = mux_in_cos477;
        10'b0111011110 : logcos3 = mux_in_cos478;
        10'b0111011111 : logcos3 = mux_in_cos479;
        10'b0111100000 : logcos3 = mux_in_cos480;
        10'b0111100001 : logcos3 = mux_in_cos481;
        10'b0111100010 : logcos3 = mux_in_cos482;
        10'b0111100011 : logcos3 = mux_in_cos483;
        10'b0111100100 : logcos3 = mux_in_cos484;
        10'b0111100101 : logcos3 = mux_in_cos485;
        10'b0111100110 : logcos3 = mux_in_cos486;
        10'b0111100111 : logcos3 = mux_in_cos487;
        10'b0111101000 : logcos3 = mux_in_cos488;
        10'b0111101001 : logcos3 = mux_in_cos489;
        10'b0111101010 : logcos3 = mux_in_cos490;
        10'b0111101011 : logcos3 = mux_in_cos491;
        10'b0111101100 : logcos3 = mux_in_cos492;
        10'b0111101101 : logcos3 = mux_in_cos493;
        10'b0111101110 : logcos3 = mux_in_cos494;
        10'b0111101111 : logcos3 = mux_in_cos495;
        10'b0111110000 : logcos3 = mux_in_cos496;
        10'b0111110001 : logcos3 = mux_in_cos497;
        10'b0111110010 : logcos3 = mux_in_cos498;
        10'b0111110011 : logcos3 = mux_in_cos499;
        10'b0111110100 : logcos3 = mux_in_cos500;
        10'b0111110101 : logcos3 = mux_in_cos501;
        10'b0111110110 : logcos3 = mux_in_cos502;
        10'b0111110111 : logcos3 = mux_in_cos503;
        10'b0111111000 : logcos3 = mux_in_cos504;
        10'b0111111001 : logcos3 = mux_in_cos505;
        10'b0111111010 : logcos3 = mux_in_cos506;
        10'b0111111011 : logcos3 = mux_in_cos507;
        10'b0111111100 : logcos3 = mux_in_cos508;
        10'b0111111101 : logcos3 = mux_in_cos509;
        10'b0111111110 : logcos3 = mux_in_cos510;
        10'b0111111111 : logcos3 = mux_in_cos511;
        10'b1000000000 : logcos3 = mux_in_cos512;
        default: logcos3 = 15'bx;
        endcase
    end

endmodule