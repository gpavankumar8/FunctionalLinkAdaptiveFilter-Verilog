`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author: Pavan Kumar
// Create Date: 29-07-2024
// Module name: log_sin_cos_LUT_8QP.v
//////////////////////////////////////////////////////////////////////////////////

module log_sin_cos_LUT_8QP
(
    input      [ 7:0] x_in1, x_in2, x_in3,
    output reg [15:0] logsin1, logsin2, logsin3, logcos1, logcos2, logcos3
);

    wire [15:0] mux_in_cos0, mux_in_sin0, mux_in_cos1, mux_in_sin1, mux_in_cos2, mux_in_sin2, mux_in_cos3, mux_in_sin3, mux_in_cos4, mux_in_sin4, mux_in_cos5, mux_in_sin5, mux_in_cos6, mux_in_sin6, mux_in_cos7, mux_in_sin7, mux_in_cos8, mux_in_sin8, mux_in_cos9, mux_in_sin9, mux_in_cos10, mux_in_sin10, mux_in_cos11, mux_in_sin11, mux_in_cos12, mux_in_sin12, mux_in_cos13, mux_in_sin13, mux_in_cos14, mux_in_sin14, mux_in_cos15, mux_in_sin15, mux_in_cos16, mux_in_sin16, mux_in_cos17, mux_in_sin17, mux_in_cos18, mux_in_sin18, mux_in_cos19, mux_in_sin19, mux_in_cos20, mux_in_sin20, mux_in_cos21, mux_in_sin21, mux_in_cos22, mux_in_sin22, mux_in_cos23, mux_in_sin23, mux_in_cos24, mux_in_sin24, mux_in_cos25, mux_in_sin25, mux_in_cos26, mux_in_sin26, mux_in_cos27, mux_in_sin27, mux_in_cos28, mux_in_sin28, mux_in_cos29, mux_in_sin29, mux_in_cos30, mux_in_sin30, mux_in_cos31, mux_in_sin31, mux_in_cos32, mux_in_sin32, mux_in_cos33, mux_in_sin33, mux_in_cos34, mux_in_sin34, mux_in_cos35, mux_in_sin35, mux_in_cos36, mux_in_sin36, mux_in_cos37, mux_in_sin37, mux_in_cos38, mux_in_sin38, mux_in_cos39, mux_in_sin39, mux_in_cos40, mux_in_sin40, mux_in_cos41, mux_in_sin41, mux_in_cos42, mux_in_sin42, mux_in_cos43, mux_in_sin43, mux_in_cos44, mux_in_sin44, mux_in_cos45, mux_in_sin45, mux_in_cos46, mux_in_sin46, mux_in_cos47, mux_in_sin47, mux_in_cos48, mux_in_sin48, mux_in_cos49, mux_in_sin49, mux_in_cos50, mux_in_sin50, mux_in_cos51, mux_in_sin51, mux_in_cos52, mux_in_sin52, mux_in_cos53, mux_in_sin53, mux_in_cos54, mux_in_sin54, mux_in_cos55, mux_in_sin55, mux_in_cos56, mux_in_sin56, mux_in_cos57, mux_in_sin57, mux_in_cos58, mux_in_sin58, mux_in_cos59, mux_in_sin59, mux_in_cos60, mux_in_sin60, mux_in_cos61, mux_in_sin61, mux_in_cos62, mux_in_sin62, mux_in_cos63, mux_in_sin63, mux_in_cos64, mux_in_sin64, mux_in_cos65, mux_in_sin65, mux_in_cos66, mux_in_sin66, mux_in_cos67, mux_in_sin67, mux_in_cos68, mux_in_sin68, mux_in_cos69, mux_in_sin69, mux_in_cos70, mux_in_sin70, mux_in_cos71, mux_in_sin71, mux_in_cos72, mux_in_sin72, mux_in_cos73, mux_in_sin73, mux_in_cos74, mux_in_sin74, mux_in_cos75, mux_in_sin75, mux_in_cos76, mux_in_sin76, mux_in_cos77, mux_in_sin77, mux_in_cos78, mux_in_sin78, mux_in_cos79, mux_in_sin79, mux_in_cos80, mux_in_sin80, mux_in_cos81, mux_in_sin81, mux_in_cos82, mux_in_sin82, mux_in_cos83, mux_in_sin83, mux_in_cos84, mux_in_sin84, mux_in_cos85, mux_in_sin85, mux_in_cos86, mux_in_sin86, mux_in_cos87, mux_in_sin87, mux_in_cos88, mux_in_sin88, mux_in_cos89, mux_in_sin89, mux_in_cos90, mux_in_sin90, mux_in_cos91, mux_in_sin91, mux_in_cos92, mux_in_sin92, mux_in_cos93, mux_in_sin93, mux_in_cos94, mux_in_sin94, mux_in_cos95, mux_in_sin95, mux_in_cos96, mux_in_sin96, mux_in_cos97, mux_in_sin97, mux_in_cos98, mux_in_sin98, mux_in_cos99, mux_in_sin99, mux_in_cos100, mux_in_sin100, mux_in_cos101, mux_in_sin101, mux_in_cos102, mux_in_sin102, mux_in_cos103, mux_in_sin103, mux_in_cos104, mux_in_sin104, mux_in_cos105, mux_in_sin105, mux_in_cos106, mux_in_sin106, mux_in_cos107, mux_in_sin107, mux_in_cos108, mux_in_sin108, mux_in_cos109, mux_in_sin109, mux_in_cos110, mux_in_sin110, mux_in_cos111, mux_in_sin111, mux_in_cos112, mux_in_sin112, mux_in_cos113, mux_in_sin113, mux_in_cos114, mux_in_sin114, mux_in_cos115, mux_in_sin115, mux_in_cos116, mux_in_sin116, mux_in_cos117, mux_in_sin117, mux_in_cos118, mux_in_sin118, mux_in_cos119, mux_in_sin119, mux_in_cos120, mux_in_sin120, mux_in_cos121, mux_in_sin121, mux_in_cos122, mux_in_sin122, mux_in_cos123, mux_in_sin123, mux_in_cos124, mux_in_sin124, mux_in_cos125, mux_in_sin125, mux_in_cos126, mux_in_sin126, mux_in_cos127, mux_in_sin127, mux_in_cos128, mux_in_sin128;

    assign mux_in_cos0 = 16'b0000000000000000;
    assign mux_in_sin0 = 16'b0000000000000000;
    assign mux_in_cos1 = 16'b0000000000000000;
    assign mux_in_sin1 = 16'b1001101001101100;
    assign mux_in_cos2 = 16'b1111111111111110;
    assign mux_in_sin2 = 16'b1010101001101100;
    assign mux_in_cos3 = 16'b1111111111111100;
    assign mux_in_sin3 = 16'b1011001111000111;
    assign mux_in_cos4 = 16'b1111111111111001;
    assign mux_in_sin4 = 16'b1011101001101010;
    assign mux_in_cos5 = 16'b1111111111110101;
    assign mux_in_sin5 = 16'b1011111110001111;
    assign mux_in_cos6 = 16'b1111111111110000;
    assign mux_in_sin6 = 16'b1100001111000011;
    assign mux_in_cos7 = 16'b1111111111101010;
    assign mux_in_sin7 = 16'b1100011101010000;
    assign mux_in_cos8 = 16'b1111111111100011;
    assign mux_in_sin8 = 16'b1100101001100011;
    assign mux_in_cos9 = 16'b1111111111011100;
    assign mux_in_sin9 = 16'b1100110100011001;
    assign mux_in_cos10 = 16'b1111111111010011;
    assign mux_in_sin10 = 16'b1100111110000100;
    assign mux_in_cos11 = 16'b1111111111001010;
    assign mux_in_sin11 = 16'b1101000110110100;
    assign mux_in_cos12 = 16'b1111111111000000;
    assign mux_in_sin12 = 16'b1101001110110011;
    assign mux_in_cos13 = 16'b1111111110110100;
    assign mux_in_sin13 = 16'b1101010110001000;
    assign mux_in_cos14 = 16'b1111111110101000;
    assign mux_in_sin14 = 16'b1101011100111010;
    assign mux_in_cos15 = 16'b1111111110011011;
    assign mux_in_sin15 = 16'b1101100011001110;
    assign mux_in_cos16 = 16'b1111111110001101;
    assign mux_in_sin16 = 16'b1101101001000111;
    assign mux_in_cos17 = 16'b1111111101111110;
    assign mux_in_sin17 = 16'b1101101110101000;
    assign mux_in_cos18 = 16'b1111111101101111;
    assign mux_in_sin18 = 16'b1101110011110100;
    assign mux_in_cos19 = 16'b1111111101011110;
    assign mux_in_sin19 = 16'b1101111000101110;
    assign mux_in_cos20 = 16'b1111111101001100;
    assign mux_in_sin20 = 16'b1101111101011000;
    assign mux_in_cos21 = 16'b1111111100111010;
    assign mux_in_sin21 = 16'b1110000001110010;
    assign mux_in_cos22 = 16'b1111111100100110;
    assign mux_in_sin22 = 16'b1110000101111110;
    assign mux_in_cos23 = 16'b1111111100010001;
    assign mux_in_sin23 = 16'b1110001001111110;
    assign mux_in_cos24 = 16'b1111111011111100;
    assign mux_in_sin24 = 16'b1110001101110011;
    assign mux_in_cos25 = 16'b1111111011100101;
    assign mux_in_sin25 = 16'b1110010001011101;
    assign mux_in_cos26 = 16'b1111111011001110;
    assign mux_in_sin26 = 16'b1110010100111101;
    assign mux_in_cos27 = 16'b1111111010110110;
    assign mux_in_sin27 = 16'b1110011000010100;
    assign mux_in_cos28 = 16'b1111111010011100;
    assign mux_in_sin28 = 16'b1110011011100011;
    assign mux_in_cos29 = 16'b1111111010000010;
    assign mux_in_sin29 = 16'b1110011110101010;
    assign mux_in_cos30 = 16'b1111111001100110;
    assign mux_in_sin30 = 16'b1110100001101001;
    assign mux_in_cos31 = 16'b1111111001001010;
    assign mux_in_sin31 = 16'b1110100100100010;
    assign mux_in_cos32 = 16'b1111111000101100;
    assign mux_in_sin32 = 16'b1110100111010100;
    assign mux_in_cos33 = 16'b1111111000001110;
    assign mux_in_sin33 = 16'b1110101010000000;
    assign mux_in_cos34 = 16'b1111110111101110;
    assign mux_in_sin34 = 16'b1110101100100110;
    assign mux_in_cos35 = 16'b1111110111001101;
    assign mux_in_sin35 = 16'b1110101111000111;
    assign mux_in_cos36 = 16'b1111110110101100;
    assign mux_in_sin36 = 16'b1110110001100011;
    assign mux_in_cos37 = 16'b1111110110001001;
    assign mux_in_sin37 = 16'b1110110011111010;
    assign mux_in_cos38 = 16'b1111110101100101;
    assign mux_in_sin38 = 16'b1110110110001100;
    assign mux_in_cos39 = 16'b1111110101000000;
    assign mux_in_sin39 = 16'b1110111000011010;
    assign mux_in_cos40 = 16'b1111110100011001;
    assign mux_in_sin40 = 16'b1110111010100100;
    assign mux_in_cos41 = 16'b1111110011110010;
    assign mux_in_sin41 = 16'b1110111100101010;
    assign mux_in_cos42 = 16'b1111110011001010;
    assign mux_in_sin42 = 16'b1110111110101011;
    assign mux_in_cos43 = 16'b1111110010100000;
    assign mux_in_sin43 = 16'b1111000000101010;
    assign mux_in_cos44 = 16'b1111110001110101;
    assign mux_in_sin44 = 16'b1111000010100100;
    assign mux_in_cos45 = 16'b1111110001001001;
    assign mux_in_sin45 = 16'b1111000100011100;
    assign mux_in_cos46 = 16'b1111110000011100;
    assign mux_in_sin46 = 16'b1111000110010000;
    assign mux_in_cos47 = 16'b1111101111101101;
    assign mux_in_sin47 = 16'b1111001000000001;
    assign mux_in_cos48 = 16'b1111101110111101;
    assign mux_in_sin48 = 16'b1111001001101111;
    assign mux_in_cos49 = 16'b1111101110001100;
    assign mux_in_sin49 = 16'b1111001011011010;
    assign mux_in_cos50 = 16'b1111101101011010;
    assign mux_in_sin50 = 16'b1111001101000010;
    assign mux_in_cos51 = 16'b1111101100100110;
    assign mux_in_sin51 = 16'b1111001110101000;
    assign mux_in_cos52 = 16'b1111101011110001;
    assign mux_in_sin52 = 16'b1111010000001011;
    assign mux_in_cos53 = 16'b1111101010111011;
    assign mux_in_sin53 = 16'b1111010001101011;
    assign mux_in_cos54 = 16'b1111101010000011;
    assign mux_in_sin54 = 16'b1111010011001010;
    assign mux_in_cos55 = 16'b1111101001001001;
    assign mux_in_sin55 = 16'b1111010100100101;
    assign mux_in_cos56 = 16'b1111101000001111;
    assign mux_in_sin56 = 16'b1111010101111111;
    assign mux_in_cos57 = 16'b1111100111010010;
    assign mux_in_sin57 = 16'b1111010111010110;
    assign mux_in_cos58 = 16'b1111100110010101;
    assign mux_in_sin58 = 16'b1111011000101011;
    assign mux_in_cos59 = 16'b1111100101010101;
    assign mux_in_sin59 = 16'b1111011001111110;
    assign mux_in_cos60 = 16'b1111100100010100;
    assign mux_in_sin60 = 16'b1111011011001111;
    assign mux_in_cos61 = 16'b1111100011010010;
    assign mux_in_sin61 = 16'b1111011100011110;
    assign mux_in_cos62 = 16'b1111100010001110;
    assign mux_in_sin62 = 16'b1111011101101011;
    assign mux_in_cos63 = 16'b1111100001001000;
    assign mux_in_sin63 = 16'b1111011110110111;
    assign mux_in_cos64 = 16'b1111100000000000;
    assign mux_in_sin64 = 16'b1111100000000000;
    assign mux_in_cos65 = 16'b1111011110110111;
    assign mux_in_sin65 = 16'b1111100001001000;
    assign mux_in_cos66 = 16'b1111011101101011;
    assign mux_in_sin66 = 16'b1111100010001110;
    assign mux_in_cos67 = 16'b1111011100011110;
    assign mux_in_sin67 = 16'b1111100011010010;
    assign mux_in_cos68 = 16'b1111011011001111;
    assign mux_in_sin68 = 16'b1111100100010100;
    assign mux_in_cos69 = 16'b1111011001111110;
    assign mux_in_sin69 = 16'b1111100101010101;
    assign mux_in_cos70 = 16'b1111011000101011;
    assign mux_in_sin70 = 16'b1111100110010101;
    assign mux_in_cos71 = 16'b1111010111010110;
    assign mux_in_sin71 = 16'b1111100111010010;
    assign mux_in_cos72 = 16'b1111010101111111;
    assign mux_in_sin72 = 16'b1111101000001111;
    assign mux_in_cos73 = 16'b1111010100100101;
    assign mux_in_sin73 = 16'b1111101001001001;
    assign mux_in_cos74 = 16'b1111010011001010;
    assign mux_in_sin74 = 16'b1111101010000011;
    assign mux_in_cos75 = 16'b1111010001101011;
    assign mux_in_sin75 = 16'b1111101010111011;
    assign mux_in_cos76 = 16'b1111010000001011;
    assign mux_in_sin76 = 16'b1111101011110001;
    assign mux_in_cos77 = 16'b1111001110101000;
    assign mux_in_sin77 = 16'b1111101100100110;
    assign mux_in_cos78 = 16'b1111001101000010;
    assign mux_in_sin78 = 16'b1111101101011010;
    assign mux_in_cos79 = 16'b1111001011011010;
    assign mux_in_sin79 = 16'b1111101110001100;
    assign mux_in_cos80 = 16'b1111001001101111;
    assign mux_in_sin80 = 16'b1111101110111101;
    assign mux_in_cos81 = 16'b1111001000000001;
    assign mux_in_sin81 = 16'b1111101111101101;
    assign mux_in_cos82 = 16'b1111000110010000;
    assign mux_in_sin82 = 16'b1111110000011100;
    assign mux_in_cos83 = 16'b1111000100011100;
    assign mux_in_sin83 = 16'b1111110001001001;
    assign mux_in_cos84 = 16'b1111000010100100;
    assign mux_in_sin84 = 16'b1111110001110101;
    assign mux_in_cos85 = 16'b1111000000101010;
    assign mux_in_sin85 = 16'b1111110010100000;
    assign mux_in_cos86 = 16'b1110111110101011;
    assign mux_in_sin86 = 16'b1111110011001010;
    assign mux_in_cos87 = 16'b1110111100101010;
    assign mux_in_sin87 = 16'b1111110011110010;
    assign mux_in_cos88 = 16'b1110111010100100;
    assign mux_in_sin88 = 16'b1111110100011001;
    assign mux_in_cos89 = 16'b1110111000011010;
    assign mux_in_sin89 = 16'b1111110101000000;
    assign mux_in_cos90 = 16'b1110110110001100;
    assign mux_in_sin90 = 16'b1111110101100101;
    assign mux_in_cos91 = 16'b1110110011111010;
    assign mux_in_sin91 = 16'b1111110110001001;
    assign mux_in_cos92 = 16'b1110110001100011;
    assign mux_in_sin92 = 16'b1111110110101100;
    assign mux_in_cos93 = 16'b1110101111000111;
    assign mux_in_sin93 = 16'b1111110111001101;
    assign mux_in_cos94 = 16'b1110101100100110;
    assign mux_in_sin94 = 16'b1111110111101110;
    assign mux_in_cos95 = 16'b1110101010000000;
    assign mux_in_sin95 = 16'b1111111000001110;
    assign mux_in_cos96 = 16'b1110100111010100;
    assign mux_in_sin96 = 16'b1111111000101100;
    assign mux_in_cos97 = 16'b1110100100100010;
    assign mux_in_sin97 = 16'b1111111001001010;
    assign mux_in_cos98 = 16'b1110100001101001;
    assign mux_in_sin98 = 16'b1111111001100110;
    assign mux_in_cos99 = 16'b1110011110101010;
    assign mux_in_sin99 = 16'b1111111010000010;
    assign mux_in_cos100 = 16'b1110011011100011;
    assign mux_in_sin100 = 16'b1111111010011100;
    assign mux_in_cos101 = 16'b1110011000010100;
    assign mux_in_sin101 = 16'b1111111010110110;
    assign mux_in_cos102 = 16'b1110010100111101;
    assign mux_in_sin102 = 16'b1111111011001110;
    assign mux_in_cos103 = 16'b1110010001011101;
    assign mux_in_sin103 = 16'b1111111011100101;
    assign mux_in_cos104 = 16'b1110001101110011;
    assign mux_in_sin104 = 16'b1111111011111100;
    assign mux_in_cos105 = 16'b1110001001111110;
    assign mux_in_sin105 = 16'b1111111100010001;
    assign mux_in_cos106 = 16'b1110000101111110;
    assign mux_in_sin106 = 16'b1111111100100110;
    assign mux_in_cos107 = 16'b1110000001110010;
    assign mux_in_sin107 = 16'b1111111100111010;
    assign mux_in_cos108 = 16'b1101111101011000;
    assign mux_in_sin108 = 16'b1111111101001100;
    assign mux_in_cos109 = 16'b1101111000101110;
    assign mux_in_sin109 = 16'b1111111101011110;
    assign mux_in_cos110 = 16'b1101110011110100;
    assign mux_in_sin110 = 16'b1111111101101111;
    assign mux_in_cos111 = 16'b1101101110101000;
    assign mux_in_sin111 = 16'b1111111101111110;
    assign mux_in_cos112 = 16'b1101101001000111;
    assign mux_in_sin112 = 16'b1111111110001101;
    assign mux_in_cos113 = 16'b1101100011001110;
    assign mux_in_sin113 = 16'b1111111110011011;
    assign mux_in_cos114 = 16'b1101011100111010;
    assign mux_in_sin114 = 16'b1111111110101000;
    assign mux_in_cos115 = 16'b1101010110001000;
    assign mux_in_sin115 = 16'b1111111110110100;
    assign mux_in_cos116 = 16'b1101001110110011;
    assign mux_in_sin116 = 16'b1111111111000000;
    assign mux_in_cos117 = 16'b1101000110110100;
    assign mux_in_sin117 = 16'b1111111111001010;
    assign mux_in_cos118 = 16'b1100111110000100;
    assign mux_in_sin118 = 16'b1111111111010011;
    assign mux_in_cos119 = 16'b1100110100011001;
    assign mux_in_sin119 = 16'b1111111111011100;
    assign mux_in_cos120 = 16'b1100101001100011;
    assign mux_in_sin120 = 16'b1111111111100011;
    assign mux_in_cos121 = 16'b1100011101010000;
    assign mux_in_sin121 = 16'b1111111111101010;
    assign mux_in_cos122 = 16'b1100001111000011;
    assign mux_in_sin122 = 16'b1111111111110000;
    assign mux_in_cos123 = 16'b1011111110001111;
    assign mux_in_sin123 = 16'b1111111111110101;
    assign mux_in_cos124 = 16'b1011101001101010;
    assign mux_in_sin124 = 16'b1111111111111001;
    assign mux_in_cos125 = 16'b1011001111000111;
    assign mux_in_sin125 = 16'b1111111111111100;
    assign mux_in_cos126 = 16'b1010101001101100;
    assign mux_in_sin126 = 16'b1111111111111110;
    assign mux_in_cos127 = 16'b1001101001101100;
    assign mux_in_sin127 = 16'b0000000000000000;
    assign mux_in_cos128 = 16'b0000000000000000;
    assign mux_in_sin128 = 16'b0000000000000000;

    always @ (*)
    begin
        case(x_in1)
        8'b00000000 : logsin1 = mux_in_sin0;
        8'b00000001 : logsin1 = mux_in_sin1;
        8'b00000010 : logsin1 = mux_in_sin2;
        8'b00000011 : logsin1 = mux_in_sin3;
        8'b00000100 : logsin1 = mux_in_sin4;
        8'b00000101 : logsin1 = mux_in_sin5;
        8'b00000110 : logsin1 = mux_in_sin6;
        8'b00000111 : logsin1 = mux_in_sin7;
        8'b00001000 : logsin1 = mux_in_sin8;
        8'b00001001 : logsin1 = mux_in_sin9;
        8'b00001010 : logsin1 = mux_in_sin10;
        8'b00001011 : logsin1 = mux_in_sin11;
        8'b00001100 : logsin1 = mux_in_sin12;
        8'b00001101 : logsin1 = mux_in_sin13;
        8'b00001110 : logsin1 = mux_in_sin14;
        8'b00001111 : logsin1 = mux_in_sin15;
        8'b00010000 : logsin1 = mux_in_sin16;
        8'b00010001 : logsin1 = mux_in_sin17;
        8'b00010010 : logsin1 = mux_in_sin18;
        8'b00010011 : logsin1 = mux_in_sin19;
        8'b00010100 : logsin1 = mux_in_sin20;
        8'b00010101 : logsin1 = mux_in_sin21;
        8'b00010110 : logsin1 = mux_in_sin22;
        8'b00010111 : logsin1 = mux_in_sin23;
        8'b00011000 : logsin1 = mux_in_sin24;
        8'b00011001 : logsin1 = mux_in_sin25;
        8'b00011010 : logsin1 = mux_in_sin26;
        8'b00011011 : logsin1 = mux_in_sin27;
        8'b00011100 : logsin1 = mux_in_sin28;
        8'b00011101 : logsin1 = mux_in_sin29;
        8'b00011110 : logsin1 = mux_in_sin30;
        8'b00011111 : logsin1 = mux_in_sin31;
        8'b00100000 : logsin1 = mux_in_sin32;
        8'b00100001 : logsin1 = mux_in_sin33;
        8'b00100010 : logsin1 = mux_in_sin34;
        8'b00100011 : logsin1 = mux_in_sin35;
        8'b00100100 : logsin1 = mux_in_sin36;
        8'b00100101 : logsin1 = mux_in_sin37;
        8'b00100110 : logsin1 = mux_in_sin38;
        8'b00100111 : logsin1 = mux_in_sin39;
        8'b00101000 : logsin1 = mux_in_sin40;
        8'b00101001 : logsin1 = mux_in_sin41;
        8'b00101010 : logsin1 = mux_in_sin42;
        8'b00101011 : logsin1 = mux_in_sin43;
        8'b00101100 : logsin1 = mux_in_sin44;
        8'b00101101 : logsin1 = mux_in_sin45;
        8'b00101110 : logsin1 = mux_in_sin46;
        8'b00101111 : logsin1 = mux_in_sin47;
        8'b00110000 : logsin1 = mux_in_sin48;
        8'b00110001 : logsin1 = mux_in_sin49;
        8'b00110010 : logsin1 = mux_in_sin50;
        8'b00110011 : logsin1 = mux_in_sin51;
        8'b00110100 : logsin1 = mux_in_sin52;
        8'b00110101 : logsin1 = mux_in_sin53;
        8'b00110110 : logsin1 = mux_in_sin54;
        8'b00110111 : logsin1 = mux_in_sin55;
        8'b00111000 : logsin1 = mux_in_sin56;
        8'b00111001 : logsin1 = mux_in_sin57;
        8'b00111010 : logsin1 = mux_in_sin58;
        8'b00111011 : logsin1 = mux_in_sin59;
        8'b00111100 : logsin1 = mux_in_sin60;
        8'b00111101 : logsin1 = mux_in_sin61;
        8'b00111110 : logsin1 = mux_in_sin62;
        8'b00111111 : logsin1 = mux_in_sin63;
        8'b01000000 : logsin1 = mux_in_sin64;
        8'b01000001 : logsin1 = mux_in_sin65;
        8'b01000010 : logsin1 = mux_in_sin66;
        8'b01000011 : logsin1 = mux_in_sin67;
        8'b01000100 : logsin1 = mux_in_sin68;
        8'b01000101 : logsin1 = mux_in_sin69;
        8'b01000110 : logsin1 = mux_in_sin70;
        8'b01000111 : logsin1 = mux_in_sin71;
        8'b01001000 : logsin1 = mux_in_sin72;
        8'b01001001 : logsin1 = mux_in_sin73;
        8'b01001010 : logsin1 = mux_in_sin74;
        8'b01001011 : logsin1 = mux_in_sin75;
        8'b01001100 : logsin1 = mux_in_sin76;
        8'b01001101 : logsin1 = mux_in_sin77;
        8'b01001110 : logsin1 = mux_in_sin78;
        8'b01001111 : logsin1 = mux_in_sin79;
        8'b01010000 : logsin1 = mux_in_sin80;
        8'b01010001 : logsin1 = mux_in_sin81;
        8'b01010010 : logsin1 = mux_in_sin82;
        8'b01010011 : logsin1 = mux_in_sin83;
        8'b01010100 : logsin1 = mux_in_sin84;
        8'b01010101 : logsin1 = mux_in_sin85;
        8'b01010110 : logsin1 = mux_in_sin86;
        8'b01010111 : logsin1 = mux_in_sin87;
        8'b01011000 : logsin1 = mux_in_sin88;
        8'b01011001 : logsin1 = mux_in_sin89;
        8'b01011010 : logsin1 = mux_in_sin90;
        8'b01011011 : logsin1 = mux_in_sin91;
        8'b01011100 : logsin1 = mux_in_sin92;
        8'b01011101 : logsin1 = mux_in_sin93;
        8'b01011110 : logsin1 = mux_in_sin94;
        8'b01011111 : logsin1 = mux_in_sin95;
        8'b01100000 : logsin1 = mux_in_sin96;
        8'b01100001 : logsin1 = mux_in_sin97;
        8'b01100010 : logsin1 = mux_in_sin98;
        8'b01100011 : logsin1 = mux_in_sin99;
        8'b01100100 : logsin1 = mux_in_sin100;
        8'b01100101 : logsin1 = mux_in_sin101;
        8'b01100110 : logsin1 = mux_in_sin102;
        8'b01100111 : logsin1 = mux_in_sin103;
        8'b01101000 : logsin1 = mux_in_sin104;
        8'b01101001 : logsin1 = mux_in_sin105;
        8'b01101010 : logsin1 = mux_in_sin106;
        8'b01101011 : logsin1 = mux_in_sin107;
        8'b01101100 : logsin1 = mux_in_sin108;
        8'b01101101 : logsin1 = mux_in_sin109;
        8'b01101110 : logsin1 = mux_in_sin110;
        8'b01101111 : logsin1 = mux_in_sin111;
        8'b01110000 : logsin1 = mux_in_sin112;
        8'b01110001 : logsin1 = mux_in_sin113;
        8'b01110010 : logsin1 = mux_in_sin114;
        8'b01110011 : logsin1 = mux_in_sin115;
        8'b01110100 : logsin1 = mux_in_sin116;
        8'b01110101 : logsin1 = mux_in_sin117;
        8'b01110110 : logsin1 = mux_in_sin118;
        8'b01110111 : logsin1 = mux_in_sin119;
        8'b01111000 : logsin1 = mux_in_sin120;
        8'b01111001 : logsin1 = mux_in_sin121;
        8'b01111010 : logsin1 = mux_in_sin122;
        8'b01111011 : logsin1 = mux_in_sin123;
        8'b01111100 : logsin1 = mux_in_sin124;
        8'b01111101 : logsin1 = mux_in_sin125;
        8'b01111110 : logsin1 = mux_in_sin126;
        8'b01111111 : logsin1 = mux_in_sin127;
        8'b10000000 : logsin1 = mux_in_sin128;
        default: logsin1 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in2)
        8'b00000000 : logsin2 = mux_in_sin0;
        8'b00000001 : logsin2 = mux_in_sin1;
        8'b00000010 : logsin2 = mux_in_sin2;
        8'b00000011 : logsin2 = mux_in_sin3;
        8'b00000100 : logsin2 = mux_in_sin4;
        8'b00000101 : logsin2 = mux_in_sin5;
        8'b00000110 : logsin2 = mux_in_sin6;
        8'b00000111 : logsin2 = mux_in_sin7;
        8'b00001000 : logsin2 = mux_in_sin8;
        8'b00001001 : logsin2 = mux_in_sin9;
        8'b00001010 : logsin2 = mux_in_sin10;
        8'b00001011 : logsin2 = mux_in_sin11;
        8'b00001100 : logsin2 = mux_in_sin12;
        8'b00001101 : logsin2 = mux_in_sin13;
        8'b00001110 : logsin2 = mux_in_sin14;
        8'b00001111 : logsin2 = mux_in_sin15;
        8'b00010000 : logsin2 = mux_in_sin16;
        8'b00010001 : logsin2 = mux_in_sin17;
        8'b00010010 : logsin2 = mux_in_sin18;
        8'b00010011 : logsin2 = mux_in_sin19;
        8'b00010100 : logsin2 = mux_in_sin20;
        8'b00010101 : logsin2 = mux_in_sin21;
        8'b00010110 : logsin2 = mux_in_sin22;
        8'b00010111 : logsin2 = mux_in_sin23;
        8'b00011000 : logsin2 = mux_in_sin24;
        8'b00011001 : logsin2 = mux_in_sin25;
        8'b00011010 : logsin2 = mux_in_sin26;
        8'b00011011 : logsin2 = mux_in_sin27;
        8'b00011100 : logsin2 = mux_in_sin28;
        8'b00011101 : logsin2 = mux_in_sin29;
        8'b00011110 : logsin2 = mux_in_sin30;
        8'b00011111 : logsin2 = mux_in_sin31;
        8'b00100000 : logsin2 = mux_in_sin32;
        8'b00100001 : logsin2 = mux_in_sin33;
        8'b00100010 : logsin2 = mux_in_sin34;
        8'b00100011 : logsin2 = mux_in_sin35;
        8'b00100100 : logsin2 = mux_in_sin36;
        8'b00100101 : logsin2 = mux_in_sin37;
        8'b00100110 : logsin2 = mux_in_sin38;
        8'b00100111 : logsin2 = mux_in_sin39;
        8'b00101000 : logsin2 = mux_in_sin40;
        8'b00101001 : logsin2 = mux_in_sin41;
        8'b00101010 : logsin2 = mux_in_sin42;
        8'b00101011 : logsin2 = mux_in_sin43;
        8'b00101100 : logsin2 = mux_in_sin44;
        8'b00101101 : logsin2 = mux_in_sin45;
        8'b00101110 : logsin2 = mux_in_sin46;
        8'b00101111 : logsin2 = mux_in_sin47;
        8'b00110000 : logsin2 = mux_in_sin48;
        8'b00110001 : logsin2 = mux_in_sin49;
        8'b00110010 : logsin2 = mux_in_sin50;
        8'b00110011 : logsin2 = mux_in_sin51;
        8'b00110100 : logsin2 = mux_in_sin52;
        8'b00110101 : logsin2 = mux_in_sin53;
        8'b00110110 : logsin2 = mux_in_sin54;
        8'b00110111 : logsin2 = mux_in_sin55;
        8'b00111000 : logsin2 = mux_in_sin56;
        8'b00111001 : logsin2 = mux_in_sin57;
        8'b00111010 : logsin2 = mux_in_sin58;
        8'b00111011 : logsin2 = mux_in_sin59;
        8'b00111100 : logsin2 = mux_in_sin60;
        8'b00111101 : logsin2 = mux_in_sin61;
        8'b00111110 : logsin2 = mux_in_sin62;
        8'b00111111 : logsin2 = mux_in_sin63;
        8'b01000000 : logsin2 = mux_in_sin64;
        8'b01000001 : logsin2 = mux_in_sin65;
        8'b01000010 : logsin2 = mux_in_sin66;
        8'b01000011 : logsin2 = mux_in_sin67;
        8'b01000100 : logsin2 = mux_in_sin68;
        8'b01000101 : logsin2 = mux_in_sin69;
        8'b01000110 : logsin2 = mux_in_sin70;
        8'b01000111 : logsin2 = mux_in_sin71;
        8'b01001000 : logsin2 = mux_in_sin72;
        8'b01001001 : logsin2 = mux_in_sin73;
        8'b01001010 : logsin2 = mux_in_sin74;
        8'b01001011 : logsin2 = mux_in_sin75;
        8'b01001100 : logsin2 = mux_in_sin76;
        8'b01001101 : logsin2 = mux_in_sin77;
        8'b01001110 : logsin2 = mux_in_sin78;
        8'b01001111 : logsin2 = mux_in_sin79;
        8'b01010000 : logsin2 = mux_in_sin80;
        8'b01010001 : logsin2 = mux_in_sin81;
        8'b01010010 : logsin2 = mux_in_sin82;
        8'b01010011 : logsin2 = mux_in_sin83;
        8'b01010100 : logsin2 = mux_in_sin84;
        8'b01010101 : logsin2 = mux_in_sin85;
        8'b01010110 : logsin2 = mux_in_sin86;
        8'b01010111 : logsin2 = mux_in_sin87;
        8'b01011000 : logsin2 = mux_in_sin88;
        8'b01011001 : logsin2 = mux_in_sin89;
        8'b01011010 : logsin2 = mux_in_sin90;
        8'b01011011 : logsin2 = mux_in_sin91;
        8'b01011100 : logsin2 = mux_in_sin92;
        8'b01011101 : logsin2 = mux_in_sin93;
        8'b01011110 : logsin2 = mux_in_sin94;
        8'b01011111 : logsin2 = mux_in_sin95;
        8'b01100000 : logsin2 = mux_in_sin96;
        8'b01100001 : logsin2 = mux_in_sin97;
        8'b01100010 : logsin2 = mux_in_sin98;
        8'b01100011 : logsin2 = mux_in_sin99;
        8'b01100100 : logsin2 = mux_in_sin100;
        8'b01100101 : logsin2 = mux_in_sin101;
        8'b01100110 : logsin2 = mux_in_sin102;
        8'b01100111 : logsin2 = mux_in_sin103;
        8'b01101000 : logsin2 = mux_in_sin104;
        8'b01101001 : logsin2 = mux_in_sin105;
        8'b01101010 : logsin2 = mux_in_sin106;
        8'b01101011 : logsin2 = mux_in_sin107;
        8'b01101100 : logsin2 = mux_in_sin108;
        8'b01101101 : logsin2 = mux_in_sin109;
        8'b01101110 : logsin2 = mux_in_sin110;
        8'b01101111 : logsin2 = mux_in_sin111;
        8'b01110000 : logsin2 = mux_in_sin112;
        8'b01110001 : logsin2 = mux_in_sin113;
        8'b01110010 : logsin2 = mux_in_sin114;
        8'b01110011 : logsin2 = mux_in_sin115;
        8'b01110100 : logsin2 = mux_in_sin116;
        8'b01110101 : logsin2 = mux_in_sin117;
        8'b01110110 : logsin2 = mux_in_sin118;
        8'b01110111 : logsin2 = mux_in_sin119;
        8'b01111000 : logsin2 = mux_in_sin120;
        8'b01111001 : logsin2 = mux_in_sin121;
        8'b01111010 : logsin2 = mux_in_sin122;
        8'b01111011 : logsin2 = mux_in_sin123;
        8'b01111100 : logsin2 = mux_in_sin124;
        8'b01111101 : logsin2 = mux_in_sin125;
        8'b01111110 : logsin2 = mux_in_sin126;
        8'b01111111 : logsin2 = mux_in_sin127;
        8'b10000000 : logsin2 = mux_in_sin128;
        default: logsin2 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in3)
        8'b00000000 : logsin3 = mux_in_sin0;
        8'b00000001 : logsin3 = mux_in_sin1;
        8'b00000010 : logsin3 = mux_in_sin2;
        8'b00000011 : logsin3 = mux_in_sin3;
        8'b00000100 : logsin3 = mux_in_sin4;
        8'b00000101 : logsin3 = mux_in_sin5;
        8'b00000110 : logsin3 = mux_in_sin6;
        8'b00000111 : logsin3 = mux_in_sin7;
        8'b00001000 : logsin3 = mux_in_sin8;
        8'b00001001 : logsin3 = mux_in_sin9;
        8'b00001010 : logsin3 = mux_in_sin10;
        8'b00001011 : logsin3 = mux_in_sin11;
        8'b00001100 : logsin3 = mux_in_sin12;
        8'b00001101 : logsin3 = mux_in_sin13;
        8'b00001110 : logsin3 = mux_in_sin14;
        8'b00001111 : logsin3 = mux_in_sin15;
        8'b00010000 : logsin3 = mux_in_sin16;
        8'b00010001 : logsin3 = mux_in_sin17;
        8'b00010010 : logsin3 = mux_in_sin18;
        8'b00010011 : logsin3 = mux_in_sin19;
        8'b00010100 : logsin3 = mux_in_sin20;
        8'b00010101 : logsin3 = mux_in_sin21;
        8'b00010110 : logsin3 = mux_in_sin22;
        8'b00010111 : logsin3 = mux_in_sin23;
        8'b00011000 : logsin3 = mux_in_sin24;
        8'b00011001 : logsin3 = mux_in_sin25;
        8'b00011010 : logsin3 = mux_in_sin26;
        8'b00011011 : logsin3 = mux_in_sin27;
        8'b00011100 : logsin3 = mux_in_sin28;
        8'b00011101 : logsin3 = mux_in_sin29;
        8'b00011110 : logsin3 = mux_in_sin30;
        8'b00011111 : logsin3 = mux_in_sin31;
        8'b00100000 : logsin3 = mux_in_sin32;
        8'b00100001 : logsin3 = mux_in_sin33;
        8'b00100010 : logsin3 = mux_in_sin34;
        8'b00100011 : logsin3 = mux_in_sin35;
        8'b00100100 : logsin3 = mux_in_sin36;
        8'b00100101 : logsin3 = mux_in_sin37;
        8'b00100110 : logsin3 = mux_in_sin38;
        8'b00100111 : logsin3 = mux_in_sin39;
        8'b00101000 : logsin3 = mux_in_sin40;
        8'b00101001 : logsin3 = mux_in_sin41;
        8'b00101010 : logsin3 = mux_in_sin42;
        8'b00101011 : logsin3 = mux_in_sin43;
        8'b00101100 : logsin3 = mux_in_sin44;
        8'b00101101 : logsin3 = mux_in_sin45;
        8'b00101110 : logsin3 = mux_in_sin46;
        8'b00101111 : logsin3 = mux_in_sin47;
        8'b00110000 : logsin3 = mux_in_sin48;
        8'b00110001 : logsin3 = mux_in_sin49;
        8'b00110010 : logsin3 = mux_in_sin50;
        8'b00110011 : logsin3 = mux_in_sin51;
        8'b00110100 : logsin3 = mux_in_sin52;
        8'b00110101 : logsin3 = mux_in_sin53;
        8'b00110110 : logsin3 = mux_in_sin54;
        8'b00110111 : logsin3 = mux_in_sin55;
        8'b00111000 : logsin3 = mux_in_sin56;
        8'b00111001 : logsin3 = mux_in_sin57;
        8'b00111010 : logsin3 = mux_in_sin58;
        8'b00111011 : logsin3 = mux_in_sin59;
        8'b00111100 : logsin3 = mux_in_sin60;
        8'b00111101 : logsin3 = mux_in_sin61;
        8'b00111110 : logsin3 = mux_in_sin62;
        8'b00111111 : logsin3 = mux_in_sin63;
        8'b01000000 : logsin3 = mux_in_sin64;
        8'b01000001 : logsin3 = mux_in_sin65;
        8'b01000010 : logsin3 = mux_in_sin66;
        8'b01000011 : logsin3 = mux_in_sin67;
        8'b01000100 : logsin3 = mux_in_sin68;
        8'b01000101 : logsin3 = mux_in_sin69;
        8'b01000110 : logsin3 = mux_in_sin70;
        8'b01000111 : logsin3 = mux_in_sin71;
        8'b01001000 : logsin3 = mux_in_sin72;
        8'b01001001 : logsin3 = mux_in_sin73;
        8'b01001010 : logsin3 = mux_in_sin74;
        8'b01001011 : logsin3 = mux_in_sin75;
        8'b01001100 : logsin3 = mux_in_sin76;
        8'b01001101 : logsin3 = mux_in_sin77;
        8'b01001110 : logsin3 = mux_in_sin78;
        8'b01001111 : logsin3 = mux_in_sin79;
        8'b01010000 : logsin3 = mux_in_sin80;
        8'b01010001 : logsin3 = mux_in_sin81;
        8'b01010010 : logsin3 = mux_in_sin82;
        8'b01010011 : logsin3 = mux_in_sin83;
        8'b01010100 : logsin3 = mux_in_sin84;
        8'b01010101 : logsin3 = mux_in_sin85;
        8'b01010110 : logsin3 = mux_in_sin86;
        8'b01010111 : logsin3 = mux_in_sin87;
        8'b01011000 : logsin3 = mux_in_sin88;
        8'b01011001 : logsin3 = mux_in_sin89;
        8'b01011010 : logsin3 = mux_in_sin90;
        8'b01011011 : logsin3 = mux_in_sin91;
        8'b01011100 : logsin3 = mux_in_sin92;
        8'b01011101 : logsin3 = mux_in_sin93;
        8'b01011110 : logsin3 = mux_in_sin94;
        8'b01011111 : logsin3 = mux_in_sin95;
        8'b01100000 : logsin3 = mux_in_sin96;
        8'b01100001 : logsin3 = mux_in_sin97;
        8'b01100010 : logsin3 = mux_in_sin98;
        8'b01100011 : logsin3 = mux_in_sin99;
        8'b01100100 : logsin3 = mux_in_sin100;
        8'b01100101 : logsin3 = mux_in_sin101;
        8'b01100110 : logsin3 = mux_in_sin102;
        8'b01100111 : logsin3 = mux_in_sin103;
        8'b01101000 : logsin3 = mux_in_sin104;
        8'b01101001 : logsin3 = mux_in_sin105;
        8'b01101010 : logsin3 = mux_in_sin106;
        8'b01101011 : logsin3 = mux_in_sin107;
        8'b01101100 : logsin3 = mux_in_sin108;
        8'b01101101 : logsin3 = mux_in_sin109;
        8'b01101110 : logsin3 = mux_in_sin110;
        8'b01101111 : logsin3 = mux_in_sin111;
        8'b01110000 : logsin3 = mux_in_sin112;
        8'b01110001 : logsin3 = mux_in_sin113;
        8'b01110010 : logsin3 = mux_in_sin114;
        8'b01110011 : logsin3 = mux_in_sin115;
        8'b01110100 : logsin3 = mux_in_sin116;
        8'b01110101 : logsin3 = mux_in_sin117;
        8'b01110110 : logsin3 = mux_in_sin118;
        8'b01110111 : logsin3 = mux_in_sin119;
        8'b01111000 : logsin3 = mux_in_sin120;
        8'b01111001 : logsin3 = mux_in_sin121;
        8'b01111010 : logsin3 = mux_in_sin122;
        8'b01111011 : logsin3 = mux_in_sin123;
        8'b01111100 : logsin3 = mux_in_sin124;
        8'b01111101 : logsin3 = mux_in_sin125;
        8'b01111110 : logsin3 = mux_in_sin126;
        8'b01111111 : logsin3 = mux_in_sin127;
        8'b10000000 : logsin3 = mux_in_sin128;
        default: logsin3 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in1)
        8'b00000000 : logcos1 = mux_in_cos0;
        8'b00000001 : logcos1 = mux_in_cos1;
        8'b00000010 : logcos1 = mux_in_cos2;
        8'b00000011 : logcos1 = mux_in_cos3;
        8'b00000100 : logcos1 = mux_in_cos4;
        8'b00000101 : logcos1 = mux_in_cos5;
        8'b00000110 : logcos1 = mux_in_cos6;
        8'b00000111 : logcos1 = mux_in_cos7;
        8'b00001000 : logcos1 = mux_in_cos8;
        8'b00001001 : logcos1 = mux_in_cos9;
        8'b00001010 : logcos1 = mux_in_cos10;
        8'b00001011 : logcos1 = mux_in_cos11;
        8'b00001100 : logcos1 = mux_in_cos12;
        8'b00001101 : logcos1 = mux_in_cos13;
        8'b00001110 : logcos1 = mux_in_cos14;
        8'b00001111 : logcos1 = mux_in_cos15;
        8'b00010000 : logcos1 = mux_in_cos16;
        8'b00010001 : logcos1 = mux_in_cos17;
        8'b00010010 : logcos1 = mux_in_cos18;
        8'b00010011 : logcos1 = mux_in_cos19;
        8'b00010100 : logcos1 = mux_in_cos20;
        8'b00010101 : logcos1 = mux_in_cos21;
        8'b00010110 : logcos1 = mux_in_cos22;
        8'b00010111 : logcos1 = mux_in_cos23;
        8'b00011000 : logcos1 = mux_in_cos24;
        8'b00011001 : logcos1 = mux_in_cos25;
        8'b00011010 : logcos1 = mux_in_cos26;
        8'b00011011 : logcos1 = mux_in_cos27;
        8'b00011100 : logcos1 = mux_in_cos28;
        8'b00011101 : logcos1 = mux_in_cos29;
        8'b00011110 : logcos1 = mux_in_cos30;
        8'b00011111 : logcos1 = mux_in_cos31;
        8'b00100000 : logcos1 = mux_in_cos32;
        8'b00100001 : logcos1 = mux_in_cos33;
        8'b00100010 : logcos1 = mux_in_cos34;
        8'b00100011 : logcos1 = mux_in_cos35;
        8'b00100100 : logcos1 = mux_in_cos36;
        8'b00100101 : logcos1 = mux_in_cos37;
        8'b00100110 : logcos1 = mux_in_cos38;
        8'b00100111 : logcos1 = mux_in_cos39;
        8'b00101000 : logcos1 = mux_in_cos40;
        8'b00101001 : logcos1 = mux_in_cos41;
        8'b00101010 : logcos1 = mux_in_cos42;
        8'b00101011 : logcos1 = mux_in_cos43;
        8'b00101100 : logcos1 = mux_in_cos44;
        8'b00101101 : logcos1 = mux_in_cos45;
        8'b00101110 : logcos1 = mux_in_cos46;
        8'b00101111 : logcos1 = mux_in_cos47;
        8'b00110000 : logcos1 = mux_in_cos48;
        8'b00110001 : logcos1 = mux_in_cos49;
        8'b00110010 : logcos1 = mux_in_cos50;
        8'b00110011 : logcos1 = mux_in_cos51;
        8'b00110100 : logcos1 = mux_in_cos52;
        8'b00110101 : logcos1 = mux_in_cos53;
        8'b00110110 : logcos1 = mux_in_cos54;
        8'b00110111 : logcos1 = mux_in_cos55;
        8'b00111000 : logcos1 = mux_in_cos56;
        8'b00111001 : logcos1 = mux_in_cos57;
        8'b00111010 : logcos1 = mux_in_cos58;
        8'b00111011 : logcos1 = mux_in_cos59;
        8'b00111100 : logcos1 = mux_in_cos60;
        8'b00111101 : logcos1 = mux_in_cos61;
        8'b00111110 : logcos1 = mux_in_cos62;
        8'b00111111 : logcos1 = mux_in_cos63;
        8'b01000000 : logcos1 = mux_in_cos64;
        8'b01000001 : logcos1 = mux_in_cos65;
        8'b01000010 : logcos1 = mux_in_cos66;
        8'b01000011 : logcos1 = mux_in_cos67;
        8'b01000100 : logcos1 = mux_in_cos68;
        8'b01000101 : logcos1 = mux_in_cos69;
        8'b01000110 : logcos1 = mux_in_cos70;
        8'b01000111 : logcos1 = mux_in_cos71;
        8'b01001000 : logcos1 = mux_in_cos72;
        8'b01001001 : logcos1 = mux_in_cos73;
        8'b01001010 : logcos1 = mux_in_cos74;
        8'b01001011 : logcos1 = mux_in_cos75;
        8'b01001100 : logcos1 = mux_in_cos76;
        8'b01001101 : logcos1 = mux_in_cos77;
        8'b01001110 : logcos1 = mux_in_cos78;
        8'b01001111 : logcos1 = mux_in_cos79;
        8'b01010000 : logcos1 = mux_in_cos80;
        8'b01010001 : logcos1 = mux_in_cos81;
        8'b01010010 : logcos1 = mux_in_cos82;
        8'b01010011 : logcos1 = mux_in_cos83;
        8'b01010100 : logcos1 = mux_in_cos84;
        8'b01010101 : logcos1 = mux_in_cos85;
        8'b01010110 : logcos1 = mux_in_cos86;
        8'b01010111 : logcos1 = mux_in_cos87;
        8'b01011000 : logcos1 = mux_in_cos88;
        8'b01011001 : logcos1 = mux_in_cos89;
        8'b01011010 : logcos1 = mux_in_cos90;
        8'b01011011 : logcos1 = mux_in_cos91;
        8'b01011100 : logcos1 = mux_in_cos92;
        8'b01011101 : logcos1 = mux_in_cos93;
        8'b01011110 : logcos1 = mux_in_cos94;
        8'b01011111 : logcos1 = mux_in_cos95;
        8'b01100000 : logcos1 = mux_in_cos96;
        8'b01100001 : logcos1 = mux_in_cos97;
        8'b01100010 : logcos1 = mux_in_cos98;
        8'b01100011 : logcos1 = mux_in_cos99;
        8'b01100100 : logcos1 = mux_in_cos100;
        8'b01100101 : logcos1 = mux_in_cos101;
        8'b01100110 : logcos1 = mux_in_cos102;
        8'b01100111 : logcos1 = mux_in_cos103;
        8'b01101000 : logcos1 = mux_in_cos104;
        8'b01101001 : logcos1 = mux_in_cos105;
        8'b01101010 : logcos1 = mux_in_cos106;
        8'b01101011 : logcos1 = mux_in_cos107;
        8'b01101100 : logcos1 = mux_in_cos108;
        8'b01101101 : logcos1 = mux_in_cos109;
        8'b01101110 : logcos1 = mux_in_cos110;
        8'b01101111 : logcos1 = mux_in_cos111;
        8'b01110000 : logcos1 = mux_in_cos112;
        8'b01110001 : logcos1 = mux_in_cos113;
        8'b01110010 : logcos1 = mux_in_cos114;
        8'b01110011 : logcos1 = mux_in_cos115;
        8'b01110100 : logcos1 = mux_in_cos116;
        8'b01110101 : logcos1 = mux_in_cos117;
        8'b01110110 : logcos1 = mux_in_cos118;
        8'b01110111 : logcos1 = mux_in_cos119;
        8'b01111000 : logcos1 = mux_in_cos120;
        8'b01111001 : logcos1 = mux_in_cos121;
        8'b01111010 : logcos1 = mux_in_cos122;
        8'b01111011 : logcos1 = mux_in_cos123;
        8'b01111100 : logcos1 = mux_in_cos124;
        8'b01111101 : logcos1 = mux_in_cos125;
        8'b01111110 : logcos1 = mux_in_cos126;
        8'b01111111 : logcos1 = mux_in_cos127;
        8'b10000000 : logcos1 = mux_in_cos128;
        default: logcos1 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in2)
        8'b00000000 : logcos2 = mux_in_cos0;
        8'b00000001 : logcos2 = mux_in_cos1;
        8'b00000010 : logcos2 = mux_in_cos2;
        8'b00000011 : logcos2 = mux_in_cos3;
        8'b00000100 : logcos2 = mux_in_cos4;
        8'b00000101 : logcos2 = mux_in_cos5;
        8'b00000110 : logcos2 = mux_in_cos6;
        8'b00000111 : logcos2 = mux_in_cos7;
        8'b00001000 : logcos2 = mux_in_cos8;
        8'b00001001 : logcos2 = mux_in_cos9;
        8'b00001010 : logcos2 = mux_in_cos10;
        8'b00001011 : logcos2 = mux_in_cos11;
        8'b00001100 : logcos2 = mux_in_cos12;
        8'b00001101 : logcos2 = mux_in_cos13;
        8'b00001110 : logcos2 = mux_in_cos14;
        8'b00001111 : logcos2 = mux_in_cos15;
        8'b00010000 : logcos2 = mux_in_cos16;
        8'b00010001 : logcos2 = mux_in_cos17;
        8'b00010010 : logcos2 = mux_in_cos18;
        8'b00010011 : logcos2 = mux_in_cos19;
        8'b00010100 : logcos2 = mux_in_cos20;
        8'b00010101 : logcos2 = mux_in_cos21;
        8'b00010110 : logcos2 = mux_in_cos22;
        8'b00010111 : logcos2 = mux_in_cos23;
        8'b00011000 : logcos2 = mux_in_cos24;
        8'b00011001 : logcos2 = mux_in_cos25;
        8'b00011010 : logcos2 = mux_in_cos26;
        8'b00011011 : logcos2 = mux_in_cos27;
        8'b00011100 : logcos2 = mux_in_cos28;
        8'b00011101 : logcos2 = mux_in_cos29;
        8'b00011110 : logcos2 = mux_in_cos30;
        8'b00011111 : logcos2 = mux_in_cos31;
        8'b00100000 : logcos2 = mux_in_cos32;
        8'b00100001 : logcos2 = mux_in_cos33;
        8'b00100010 : logcos2 = mux_in_cos34;
        8'b00100011 : logcos2 = mux_in_cos35;
        8'b00100100 : logcos2 = mux_in_cos36;
        8'b00100101 : logcos2 = mux_in_cos37;
        8'b00100110 : logcos2 = mux_in_cos38;
        8'b00100111 : logcos2 = mux_in_cos39;
        8'b00101000 : logcos2 = mux_in_cos40;
        8'b00101001 : logcos2 = mux_in_cos41;
        8'b00101010 : logcos2 = mux_in_cos42;
        8'b00101011 : logcos2 = mux_in_cos43;
        8'b00101100 : logcos2 = mux_in_cos44;
        8'b00101101 : logcos2 = mux_in_cos45;
        8'b00101110 : logcos2 = mux_in_cos46;
        8'b00101111 : logcos2 = mux_in_cos47;
        8'b00110000 : logcos2 = mux_in_cos48;
        8'b00110001 : logcos2 = mux_in_cos49;
        8'b00110010 : logcos2 = mux_in_cos50;
        8'b00110011 : logcos2 = mux_in_cos51;
        8'b00110100 : logcos2 = mux_in_cos52;
        8'b00110101 : logcos2 = mux_in_cos53;
        8'b00110110 : logcos2 = mux_in_cos54;
        8'b00110111 : logcos2 = mux_in_cos55;
        8'b00111000 : logcos2 = mux_in_cos56;
        8'b00111001 : logcos2 = mux_in_cos57;
        8'b00111010 : logcos2 = mux_in_cos58;
        8'b00111011 : logcos2 = mux_in_cos59;
        8'b00111100 : logcos2 = mux_in_cos60;
        8'b00111101 : logcos2 = mux_in_cos61;
        8'b00111110 : logcos2 = mux_in_cos62;
        8'b00111111 : logcos2 = mux_in_cos63;
        8'b01000000 : logcos2 = mux_in_cos64;
        8'b01000001 : logcos2 = mux_in_cos65;
        8'b01000010 : logcos2 = mux_in_cos66;
        8'b01000011 : logcos2 = mux_in_cos67;
        8'b01000100 : logcos2 = mux_in_cos68;
        8'b01000101 : logcos2 = mux_in_cos69;
        8'b01000110 : logcos2 = mux_in_cos70;
        8'b01000111 : logcos2 = mux_in_cos71;
        8'b01001000 : logcos2 = mux_in_cos72;
        8'b01001001 : logcos2 = mux_in_cos73;
        8'b01001010 : logcos2 = mux_in_cos74;
        8'b01001011 : logcos2 = mux_in_cos75;
        8'b01001100 : logcos2 = mux_in_cos76;
        8'b01001101 : logcos2 = mux_in_cos77;
        8'b01001110 : logcos2 = mux_in_cos78;
        8'b01001111 : logcos2 = mux_in_cos79;
        8'b01010000 : logcos2 = mux_in_cos80;
        8'b01010001 : logcos2 = mux_in_cos81;
        8'b01010010 : logcos2 = mux_in_cos82;
        8'b01010011 : logcos2 = mux_in_cos83;
        8'b01010100 : logcos2 = mux_in_cos84;
        8'b01010101 : logcos2 = mux_in_cos85;
        8'b01010110 : logcos2 = mux_in_cos86;
        8'b01010111 : logcos2 = mux_in_cos87;
        8'b01011000 : logcos2 = mux_in_cos88;
        8'b01011001 : logcos2 = mux_in_cos89;
        8'b01011010 : logcos2 = mux_in_cos90;
        8'b01011011 : logcos2 = mux_in_cos91;
        8'b01011100 : logcos2 = mux_in_cos92;
        8'b01011101 : logcos2 = mux_in_cos93;
        8'b01011110 : logcos2 = mux_in_cos94;
        8'b01011111 : logcos2 = mux_in_cos95;
        8'b01100000 : logcos2 = mux_in_cos96;
        8'b01100001 : logcos2 = mux_in_cos97;
        8'b01100010 : logcos2 = mux_in_cos98;
        8'b01100011 : logcos2 = mux_in_cos99;
        8'b01100100 : logcos2 = mux_in_cos100;
        8'b01100101 : logcos2 = mux_in_cos101;
        8'b01100110 : logcos2 = mux_in_cos102;
        8'b01100111 : logcos2 = mux_in_cos103;
        8'b01101000 : logcos2 = mux_in_cos104;
        8'b01101001 : logcos2 = mux_in_cos105;
        8'b01101010 : logcos2 = mux_in_cos106;
        8'b01101011 : logcos2 = mux_in_cos107;
        8'b01101100 : logcos2 = mux_in_cos108;
        8'b01101101 : logcos2 = mux_in_cos109;
        8'b01101110 : logcos2 = mux_in_cos110;
        8'b01101111 : logcos2 = mux_in_cos111;
        8'b01110000 : logcos2 = mux_in_cos112;
        8'b01110001 : logcos2 = mux_in_cos113;
        8'b01110010 : logcos2 = mux_in_cos114;
        8'b01110011 : logcos2 = mux_in_cos115;
        8'b01110100 : logcos2 = mux_in_cos116;
        8'b01110101 : logcos2 = mux_in_cos117;
        8'b01110110 : logcos2 = mux_in_cos118;
        8'b01110111 : logcos2 = mux_in_cos119;
        8'b01111000 : logcos2 = mux_in_cos120;
        8'b01111001 : logcos2 = mux_in_cos121;
        8'b01111010 : logcos2 = mux_in_cos122;
        8'b01111011 : logcos2 = mux_in_cos123;
        8'b01111100 : logcos2 = mux_in_cos124;
        8'b01111101 : logcos2 = mux_in_cos125;
        8'b01111110 : logcos2 = mux_in_cos126;
        8'b01111111 : logcos2 = mux_in_cos127;
        8'b10000000 : logcos2 = mux_in_cos128;
        default: logcos2 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in3)
        8'b00000000 : logcos3 = mux_in_cos0;
        8'b00000001 : logcos3 = mux_in_cos1;
        8'b00000010 : logcos3 = mux_in_cos2;
        8'b00000011 : logcos3 = mux_in_cos3;
        8'b00000100 : logcos3 = mux_in_cos4;
        8'b00000101 : logcos3 = mux_in_cos5;
        8'b00000110 : logcos3 = mux_in_cos6;
        8'b00000111 : logcos3 = mux_in_cos7;
        8'b00001000 : logcos3 = mux_in_cos8;
        8'b00001001 : logcos3 = mux_in_cos9;
        8'b00001010 : logcos3 = mux_in_cos10;
        8'b00001011 : logcos3 = mux_in_cos11;
        8'b00001100 : logcos3 = mux_in_cos12;
        8'b00001101 : logcos3 = mux_in_cos13;
        8'b00001110 : logcos3 = mux_in_cos14;
        8'b00001111 : logcos3 = mux_in_cos15;
        8'b00010000 : logcos3 = mux_in_cos16;
        8'b00010001 : logcos3 = mux_in_cos17;
        8'b00010010 : logcos3 = mux_in_cos18;
        8'b00010011 : logcos3 = mux_in_cos19;
        8'b00010100 : logcos3 = mux_in_cos20;
        8'b00010101 : logcos3 = mux_in_cos21;
        8'b00010110 : logcos3 = mux_in_cos22;
        8'b00010111 : logcos3 = mux_in_cos23;
        8'b00011000 : logcos3 = mux_in_cos24;
        8'b00011001 : logcos3 = mux_in_cos25;
        8'b00011010 : logcos3 = mux_in_cos26;
        8'b00011011 : logcos3 = mux_in_cos27;
        8'b00011100 : logcos3 = mux_in_cos28;
        8'b00011101 : logcos3 = mux_in_cos29;
        8'b00011110 : logcos3 = mux_in_cos30;
        8'b00011111 : logcos3 = mux_in_cos31;
        8'b00100000 : logcos3 = mux_in_cos32;
        8'b00100001 : logcos3 = mux_in_cos33;
        8'b00100010 : logcos3 = mux_in_cos34;
        8'b00100011 : logcos3 = mux_in_cos35;
        8'b00100100 : logcos3 = mux_in_cos36;
        8'b00100101 : logcos3 = mux_in_cos37;
        8'b00100110 : logcos3 = mux_in_cos38;
        8'b00100111 : logcos3 = mux_in_cos39;
        8'b00101000 : logcos3 = mux_in_cos40;
        8'b00101001 : logcos3 = mux_in_cos41;
        8'b00101010 : logcos3 = mux_in_cos42;
        8'b00101011 : logcos3 = mux_in_cos43;
        8'b00101100 : logcos3 = mux_in_cos44;
        8'b00101101 : logcos3 = mux_in_cos45;
        8'b00101110 : logcos3 = mux_in_cos46;
        8'b00101111 : logcos3 = mux_in_cos47;
        8'b00110000 : logcos3 = mux_in_cos48;
        8'b00110001 : logcos3 = mux_in_cos49;
        8'b00110010 : logcos3 = mux_in_cos50;
        8'b00110011 : logcos3 = mux_in_cos51;
        8'b00110100 : logcos3 = mux_in_cos52;
        8'b00110101 : logcos3 = mux_in_cos53;
        8'b00110110 : logcos3 = mux_in_cos54;
        8'b00110111 : logcos3 = mux_in_cos55;
        8'b00111000 : logcos3 = mux_in_cos56;
        8'b00111001 : logcos3 = mux_in_cos57;
        8'b00111010 : logcos3 = mux_in_cos58;
        8'b00111011 : logcos3 = mux_in_cos59;
        8'b00111100 : logcos3 = mux_in_cos60;
        8'b00111101 : logcos3 = mux_in_cos61;
        8'b00111110 : logcos3 = mux_in_cos62;
        8'b00111111 : logcos3 = mux_in_cos63;
        8'b01000000 : logcos3 = mux_in_cos64;
        8'b01000001 : logcos3 = mux_in_cos65;
        8'b01000010 : logcos3 = mux_in_cos66;
        8'b01000011 : logcos3 = mux_in_cos67;
        8'b01000100 : logcos3 = mux_in_cos68;
        8'b01000101 : logcos3 = mux_in_cos69;
        8'b01000110 : logcos3 = mux_in_cos70;
        8'b01000111 : logcos3 = mux_in_cos71;
        8'b01001000 : logcos3 = mux_in_cos72;
        8'b01001001 : logcos3 = mux_in_cos73;
        8'b01001010 : logcos3 = mux_in_cos74;
        8'b01001011 : logcos3 = mux_in_cos75;
        8'b01001100 : logcos3 = mux_in_cos76;
        8'b01001101 : logcos3 = mux_in_cos77;
        8'b01001110 : logcos3 = mux_in_cos78;
        8'b01001111 : logcos3 = mux_in_cos79;
        8'b01010000 : logcos3 = mux_in_cos80;
        8'b01010001 : logcos3 = mux_in_cos81;
        8'b01010010 : logcos3 = mux_in_cos82;
        8'b01010011 : logcos3 = mux_in_cos83;
        8'b01010100 : logcos3 = mux_in_cos84;
        8'b01010101 : logcos3 = mux_in_cos85;
        8'b01010110 : logcos3 = mux_in_cos86;
        8'b01010111 : logcos3 = mux_in_cos87;
        8'b01011000 : logcos3 = mux_in_cos88;
        8'b01011001 : logcos3 = mux_in_cos89;
        8'b01011010 : logcos3 = mux_in_cos90;
        8'b01011011 : logcos3 = mux_in_cos91;
        8'b01011100 : logcos3 = mux_in_cos92;
        8'b01011101 : logcos3 = mux_in_cos93;
        8'b01011110 : logcos3 = mux_in_cos94;
        8'b01011111 : logcos3 = mux_in_cos95;
        8'b01100000 : logcos3 = mux_in_cos96;
        8'b01100001 : logcos3 = mux_in_cos97;
        8'b01100010 : logcos3 = mux_in_cos98;
        8'b01100011 : logcos3 = mux_in_cos99;
        8'b01100100 : logcos3 = mux_in_cos100;
        8'b01100101 : logcos3 = mux_in_cos101;
        8'b01100110 : logcos3 = mux_in_cos102;
        8'b01100111 : logcos3 = mux_in_cos103;
        8'b01101000 : logcos3 = mux_in_cos104;
        8'b01101001 : logcos3 = mux_in_cos105;
        8'b01101010 : logcos3 = mux_in_cos106;
        8'b01101011 : logcos3 = mux_in_cos107;
        8'b01101100 : logcos3 = mux_in_cos108;
        8'b01101101 : logcos3 = mux_in_cos109;
        8'b01101110 : logcos3 = mux_in_cos110;
        8'b01101111 : logcos3 = mux_in_cos111;
        8'b01110000 : logcos3 = mux_in_cos112;
        8'b01110001 : logcos3 = mux_in_cos113;
        8'b01110010 : logcos3 = mux_in_cos114;
        8'b01110011 : logcos3 = mux_in_cos115;
        8'b01110100 : logcos3 = mux_in_cos116;
        8'b01110101 : logcos3 = mux_in_cos117;
        8'b01110110 : logcos3 = mux_in_cos118;
        8'b01110111 : logcos3 = mux_in_cos119;
        8'b01111000 : logcos3 = mux_in_cos120;
        8'b01111001 : logcos3 = mux_in_cos121;
        8'b01111010 : logcos3 = mux_in_cos122;
        8'b01111011 : logcos3 = mux_in_cos123;
        8'b01111100 : logcos3 = mux_in_cos124;
        8'b01111101 : logcos3 = mux_in_cos125;
        8'b01111110 : logcos3 = mux_in_cos126;
        8'b01111111 : logcos3 = mux_in_cos127;
        8'b10000000 : logcos3 = mux_in_cos128;
        default: logcos3 = 15'bx;
        endcase
    end
    
endmodule