`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author: Pavan Kumar
// Create Date: 10-07-2022
// Module name: sin_cos_LUT_8QP.v
//////////////////////////////////////////////////////////////////////////////////

module sin_cos_LUT_8QP
(
    input      [ 7:0] x_in1, x_in2, x_in3,
    output reg [15:0] sin1, sin2, sin3, cos1, cos2, cos3
);

    wire [15:0] mux_in_cos0, mux_in_sin0, mux_in_cos1, mux_in_sin1, mux_in_cos2, mux_in_sin2, mux_in_cos3, mux_in_sin3, mux_in_cos4, mux_in_sin4, mux_in_cos5, mux_in_sin5, mux_in_cos6, mux_in_sin6, mux_in_cos7, mux_in_sin7, mux_in_cos8, mux_in_sin8, mux_in_cos9, mux_in_sin9, mux_in_cos10, mux_in_sin10, mux_in_cos11, mux_in_sin11, mux_in_cos12, mux_in_sin12, mux_in_cos13, mux_in_sin13, mux_in_cos14, mux_in_sin14, mux_in_cos15, mux_in_sin15, mux_in_cos16, mux_in_sin16, mux_in_cos17, mux_in_sin17, mux_in_cos18, mux_in_sin18, mux_in_cos19, mux_in_sin19, mux_in_cos20, mux_in_sin20, mux_in_cos21, mux_in_sin21, mux_in_cos22, mux_in_sin22, mux_in_cos23, mux_in_sin23, mux_in_cos24, mux_in_sin24, mux_in_cos25, mux_in_sin25, mux_in_cos26, mux_in_sin26, mux_in_cos27, mux_in_sin27, mux_in_cos28, mux_in_sin28, mux_in_cos29, mux_in_sin29, mux_in_cos30, mux_in_sin30, mux_in_cos31, mux_in_sin31, mux_in_cos32, mux_in_sin32, mux_in_cos33, mux_in_sin33, mux_in_cos34, mux_in_sin34, mux_in_cos35, mux_in_sin35, mux_in_cos36, mux_in_sin36, mux_in_cos37, mux_in_sin37, mux_in_cos38, mux_in_sin38, mux_in_cos39, mux_in_sin39, mux_in_cos40, mux_in_sin40, mux_in_cos41, mux_in_sin41, mux_in_cos42, mux_in_sin42, mux_in_cos43, mux_in_sin43, mux_in_cos44, mux_in_sin44, mux_in_cos45, mux_in_sin45, mux_in_cos46, mux_in_sin46, mux_in_cos47, mux_in_sin47, mux_in_cos48, mux_in_sin48, mux_in_cos49, mux_in_sin49, mux_in_cos50, mux_in_sin50, mux_in_cos51, mux_in_sin51, mux_in_cos52, mux_in_sin52, mux_in_cos53, mux_in_sin53, mux_in_cos54, mux_in_sin54, mux_in_cos55, mux_in_sin55, mux_in_cos56, mux_in_sin56, mux_in_cos57, mux_in_sin57, mux_in_cos58, mux_in_sin58, mux_in_cos59, mux_in_sin59, mux_in_cos60, mux_in_sin60, mux_in_cos61, mux_in_sin61, mux_in_cos62, mux_in_sin62, mux_in_cos63, mux_in_sin63, mux_in_cos64, mux_in_sin64, mux_in_cos65, mux_in_sin65, mux_in_cos66, mux_in_sin66, mux_in_cos67, mux_in_sin67, mux_in_cos68, mux_in_sin68, mux_in_cos69, mux_in_sin69, mux_in_cos70, mux_in_sin70, mux_in_cos71, mux_in_sin71, mux_in_cos72, mux_in_sin72, mux_in_cos73, mux_in_sin73, mux_in_cos74, mux_in_sin74, mux_in_cos75, mux_in_sin75, mux_in_cos76, mux_in_sin76, mux_in_cos77, mux_in_sin77, mux_in_cos78, mux_in_sin78, mux_in_cos79, mux_in_sin79, mux_in_cos80, mux_in_sin80, mux_in_cos81, mux_in_sin81, mux_in_cos82, mux_in_sin82, mux_in_cos83, mux_in_sin83, mux_in_cos84, mux_in_sin84, mux_in_cos85, mux_in_sin85, mux_in_cos86, mux_in_sin86, mux_in_cos87, mux_in_sin87, mux_in_cos88, mux_in_sin88, mux_in_cos89, mux_in_sin89, mux_in_cos90, mux_in_sin90, mux_in_cos91, mux_in_sin91, mux_in_cos92, mux_in_sin92, mux_in_cos93, mux_in_sin93, mux_in_cos94, mux_in_sin94, mux_in_cos95, mux_in_sin95, mux_in_cos96, mux_in_sin96, mux_in_cos97, mux_in_sin97, mux_in_cos98, mux_in_sin98, mux_in_cos99, mux_in_sin99, mux_in_cos100, mux_in_sin100, mux_in_cos101, mux_in_sin101, mux_in_cos102, mux_in_sin102, mux_in_cos103, mux_in_sin103, mux_in_cos104, mux_in_sin104, mux_in_cos105, mux_in_sin105, mux_in_cos106, mux_in_sin106, mux_in_cos107, mux_in_sin107, mux_in_cos108, mux_in_sin108, mux_in_cos109, mux_in_sin109, mux_in_cos110, mux_in_sin110, mux_in_cos111, mux_in_sin111, mux_in_cos112, mux_in_sin112, mux_in_cos113, mux_in_sin113, mux_in_cos114, mux_in_sin114, mux_in_cos115, mux_in_sin115, mux_in_cos116, mux_in_sin116, mux_in_cos117, mux_in_sin117, mux_in_cos118, mux_in_sin118, mux_in_cos119, mux_in_sin119, mux_in_cos120, mux_in_sin120, mux_in_cos121, mux_in_sin121, mux_in_cos122, mux_in_sin122, mux_in_cos123, mux_in_sin123, mux_in_cos124, mux_in_sin124, mux_in_cos125, mux_in_sin125, mux_in_cos126, mux_in_sin126, mux_in_cos127, mux_in_sin127, mux_in_cos128, mux_in_sin128;

    assign mux_in_cos0 = 16'b1000000000000000;
    assign mux_in_sin0 = 16'b0000000000000000;
    assign mux_in_cos1 = 16'b0111111111111110;
    assign mux_in_sin1 = 16'b0000000110010010;
    assign mux_in_cos2 = 16'b0111111111110110;
    assign mux_in_sin2 = 16'b0000001100100100;
    assign mux_in_cos3 = 16'b0111111111101010;
    assign mux_in_sin3 = 16'b0000010010110110;
    assign mux_in_cos4 = 16'b0111111111011001;
    assign mux_in_sin4 = 16'b0000011001001000;
    assign mux_in_cos5 = 16'b0111111111000010;
    assign mux_in_sin5 = 16'b0000011111011001;
    assign mux_in_cos6 = 16'b0111111110100111;
    assign mux_in_sin6 = 16'b0000100101101011;
    assign mux_in_cos7 = 16'b0111111110000111;
    assign mux_in_sin7 = 16'b0000101011111011;
    assign mux_in_cos8 = 16'b0111111101100010;
    assign mux_in_sin8 = 16'b0000110010001100;
    assign mux_in_cos9 = 16'b0111111100111000;
    assign mux_in_sin9 = 16'b0000111000011100;
    assign mux_in_cos10 = 16'b0111111100001010;
    assign mux_in_sin10 = 16'b0000111110101011;
    assign mux_in_cos11 = 16'b0111111011010110;
    assign mux_in_sin11 = 16'b0001000100111010;
    assign mux_in_cos12 = 16'b0111111010011101;
    assign mux_in_sin12 = 16'b0001001011001000;
    assign mux_in_cos13 = 16'b0111111001100000;
    assign mux_in_sin13 = 16'b0001010001010101;
    assign mux_in_cos14 = 16'b0111111000011110;
    assign mux_in_sin14 = 16'b0001010111100010;
    assign mux_in_cos15 = 16'b0111110111010110;
    assign mux_in_sin15 = 16'b0001011101101110;
    assign mux_in_cos16 = 16'b0111110110001010;
    assign mux_in_sin16 = 16'b0001100011111001;
    assign mux_in_cos17 = 16'b0111110100111010;
    assign mux_in_sin17 = 16'b0001101010000011;
    assign mux_in_cos18 = 16'b0111110011100100;
    assign mux_in_sin18 = 16'b0001110000001100;
    assign mux_in_cos19 = 16'b0111110010001001;
    assign mux_in_sin19 = 16'b0001110110010011;
    assign mux_in_cos20 = 16'b0111110000101010;
    assign mux_in_sin20 = 16'b0001111100011010;
    assign mux_in_cos21 = 16'b0111101111000110;
    assign mux_in_sin21 = 16'b0010000010011111;
    assign mux_in_cos22 = 16'b0111101101011101;
    assign mux_in_sin22 = 16'b0010001000100100;
    assign mux_in_cos23 = 16'b0111101011101111;
    assign mux_in_sin23 = 16'b0010001110100111;
    assign mux_in_cos24 = 16'b0111101001111101;
    assign mux_in_sin24 = 16'b0010010100101000;
    assign mux_in_cos25 = 16'b0111101000000110;
    assign mux_in_sin25 = 16'b0010011010101000;
    assign mux_in_cos26 = 16'b0111100110001010;
    assign mux_in_sin26 = 16'b0010100000100111;
    assign mux_in_cos27 = 16'b0111100100001010;
    assign mux_in_sin27 = 16'b0010100110100100;
    assign mux_in_cos28 = 16'b0111100010000101;
    assign mux_in_sin28 = 16'b0010101100011111;
    assign mux_in_cos29 = 16'b0111011111111011;
    assign mux_in_sin29 = 16'b0010110010011001;
    assign mux_in_cos30 = 16'b0111011101101100;
    assign mux_in_sin30 = 16'b0010111000010001;
    assign mux_in_cos31 = 16'b0111011011011001;
    assign mux_in_sin31 = 16'b0010111110000111;
    assign mux_in_cos32 = 16'b0111011001000010;
    assign mux_in_sin32 = 16'b0011000011111100;
    assign mux_in_cos33 = 16'b0111010110100110;
    assign mux_in_sin33 = 16'b0011001001101110;
    assign mux_in_cos34 = 16'b0111010100000101;
    assign mux_in_sin34 = 16'b0011001111011111;
    assign mux_in_cos35 = 16'b0111010001100000;
    assign mux_in_sin35 = 16'b0011010101001110;
    assign mux_in_cos36 = 16'b0111001110110110;
    assign mux_in_sin36 = 16'b0011011010111010;
    assign mux_in_cos37 = 16'b0111001100001000;
    assign mux_in_sin37 = 16'b0011100000100101;
    assign mux_in_cos38 = 16'b0111001001010101;
    assign mux_in_sin38 = 16'b0011100110001101;
    assign mux_in_cos39 = 16'b0111000110011110;
    assign mux_in_sin39 = 16'b0011101011110011;
    assign mux_in_cos40 = 16'b0111000011100011;
    assign mux_in_sin40 = 16'b0011110001010111;
    assign mux_in_cos41 = 16'b0111000000100011;
    assign mux_in_sin41 = 16'b0011110110111000;
    assign mux_in_cos42 = 16'b0110111101011111;
    assign mux_in_sin42 = 16'b0011111100010111;
    assign mux_in_cos43 = 16'b0110111010010111;
    assign mux_in_sin43 = 16'b0100000001110100;
    assign mux_in_cos44 = 16'b0110110111001010;
    assign mux_in_sin44 = 16'b0100000111001110;
    assign mux_in_cos45 = 16'b0110110011111001;
    assign mux_in_sin45 = 16'b0100001100100110;
    assign mux_in_cos46 = 16'b0110110000100100;
    assign mux_in_sin46 = 16'b0100010001111011;
    assign mux_in_cos47 = 16'b0110101101001011;
    assign mux_in_sin47 = 16'b0100010111001101;
    assign mux_in_cos48 = 16'b0110101001101110;
    assign mux_in_sin48 = 16'b0100011100011101;
    assign mux_in_cos49 = 16'b0110100110001100;
    assign mux_in_sin49 = 16'b0100100001101010;
    assign mux_in_cos50 = 16'b0110100010100111;
    assign mux_in_sin50 = 16'b0100100110110100;
    assign mux_in_cos51 = 16'b0110011110111101;
    assign mux_in_sin51 = 16'b0100101011111011;
    assign mux_in_cos52 = 16'b0110011011010000;
    assign mux_in_sin52 = 16'b0100110001000000;
    assign mux_in_cos53 = 16'b0110010111011110;
    assign mux_in_sin53 = 16'b0100110110000001;
    assign mux_in_cos54 = 16'b0110010011101001;
    assign mux_in_sin54 = 16'b0100111011000000;
    assign mux_in_cos55 = 16'b0110001111101111;
    assign mux_in_sin55 = 16'b0100111111111011;
    assign mux_in_cos56 = 16'b0110001011110010;
    assign mux_in_sin56 = 16'b0101000100110100;
    assign mux_in_cos57 = 16'b0110000111110001;
    assign mux_in_sin57 = 16'b0101001001101001;
    assign mux_in_cos58 = 16'b0110000011101100;
    assign mux_in_sin58 = 16'b0101001110011011;
    assign mux_in_cos59 = 16'b0101111111100100;
    assign mux_in_sin59 = 16'b0101010011001010;
    assign mux_in_cos60 = 16'b0101111011010111;
    assign mux_in_sin60 = 16'b0101010111110110;
    assign mux_in_cos61 = 16'b0101110111001000;
    assign mux_in_sin61 = 16'b0101011100011110;
    assign mux_in_cos62 = 16'b0101110010110100;
    assign mux_in_sin62 = 16'b0101100001000011;
    assign mux_in_cos63 = 16'b0101101110011101;
    assign mux_in_sin63 = 16'b0101100101100100;
    assign mux_in_cos64 = 16'b0101101010000010;
    assign mux_in_sin64 = 16'b0101101010000010;
    assign mux_in_cos65 = 16'b0101100101100100;
    assign mux_in_sin65 = 16'b0101101110011101;
    assign mux_in_cos66 = 16'b0101100001000011;
    assign mux_in_sin66 = 16'b0101110010110100;
    assign mux_in_cos67 = 16'b0101011100011110;
    assign mux_in_sin67 = 16'b0101110111001000;
    assign mux_in_cos68 = 16'b0101010111110110;
    assign mux_in_sin68 = 16'b0101111011010111;
    assign mux_in_cos69 = 16'b0101010011001010;
    assign mux_in_sin69 = 16'b0101111111100100;
    assign mux_in_cos70 = 16'b0101001110011011;
    assign mux_in_sin70 = 16'b0110000011101100;
    assign mux_in_cos71 = 16'b0101001001101001;
    assign mux_in_sin71 = 16'b0110000111110001;
    assign mux_in_cos72 = 16'b0101000100110100;
    assign mux_in_sin72 = 16'b0110001011110010;
    assign mux_in_cos73 = 16'b0100111111111011;
    assign mux_in_sin73 = 16'b0110001111101111;
    assign mux_in_cos74 = 16'b0100111011000000;
    assign mux_in_sin74 = 16'b0110010011101001;
    assign mux_in_cos75 = 16'b0100110110000001;
    assign mux_in_sin75 = 16'b0110010111011110;
    assign mux_in_cos76 = 16'b0100110001000000;
    assign mux_in_sin76 = 16'b0110011011010000;
    assign mux_in_cos77 = 16'b0100101011111011;
    assign mux_in_sin77 = 16'b0110011110111101;
    assign mux_in_cos78 = 16'b0100100110110100;
    assign mux_in_sin78 = 16'b0110100010100111;
    assign mux_in_cos79 = 16'b0100100001101010;
    assign mux_in_sin79 = 16'b0110100110001100;
    assign mux_in_cos80 = 16'b0100011100011101;
    assign mux_in_sin80 = 16'b0110101001101110;
    assign mux_in_cos81 = 16'b0100010111001101;
    assign mux_in_sin81 = 16'b0110101101001011;
    assign mux_in_cos82 = 16'b0100010001111011;
    assign mux_in_sin82 = 16'b0110110000100100;
    assign mux_in_cos83 = 16'b0100001100100110;
    assign mux_in_sin83 = 16'b0110110011111001;
    assign mux_in_cos84 = 16'b0100000111001110;
    assign mux_in_sin84 = 16'b0110110111001010;
    assign mux_in_cos85 = 16'b0100000001110100;
    assign mux_in_sin85 = 16'b0110111010010111;
    assign mux_in_cos86 = 16'b0011111100010111;
    assign mux_in_sin86 = 16'b0110111101011111;
    assign mux_in_cos87 = 16'b0011110110111000;
    assign mux_in_sin87 = 16'b0111000000100011;
    assign mux_in_cos88 = 16'b0011110001010111;
    assign mux_in_sin88 = 16'b0111000011100011;
    assign mux_in_cos89 = 16'b0011101011110011;
    assign mux_in_sin89 = 16'b0111000110011110;
    assign mux_in_cos90 = 16'b0011100110001101;
    assign mux_in_sin90 = 16'b0111001001010101;
    assign mux_in_cos91 = 16'b0011100000100101;
    assign mux_in_sin91 = 16'b0111001100001000;
    assign mux_in_cos92 = 16'b0011011010111010;
    assign mux_in_sin92 = 16'b0111001110110110;
    assign mux_in_cos93 = 16'b0011010101001110;
    assign mux_in_sin93 = 16'b0111010001100000;
    assign mux_in_cos94 = 16'b0011001111011111;
    assign mux_in_sin94 = 16'b0111010100000101;
    assign mux_in_cos95 = 16'b0011001001101110;
    assign mux_in_sin95 = 16'b0111010110100110;
    assign mux_in_cos96 = 16'b0011000011111100;
    assign mux_in_sin96 = 16'b0111011001000010;
    assign mux_in_cos97 = 16'b0010111110000111;
    assign mux_in_sin97 = 16'b0111011011011001;
    assign mux_in_cos98 = 16'b0010111000010001;
    assign mux_in_sin98 = 16'b0111011101101100;
    assign mux_in_cos99 = 16'b0010110010011001;
    assign mux_in_sin99 = 16'b0111011111111011;
    assign mux_in_cos100 = 16'b0010101100011111;
    assign mux_in_sin100 = 16'b0111100010000101;
    assign mux_in_cos101 = 16'b0010100110100100;
    assign mux_in_sin101 = 16'b0111100100001010;
    assign mux_in_cos102 = 16'b0010100000100111;
    assign mux_in_sin102 = 16'b0111100110001010;
    assign mux_in_cos103 = 16'b0010011010101000;
    assign mux_in_sin103 = 16'b0111101000000110;
    assign mux_in_cos104 = 16'b0010010100101000;
    assign mux_in_sin104 = 16'b0111101001111101;
    assign mux_in_cos105 = 16'b0010001110100111;
    assign mux_in_sin105 = 16'b0111101011101111;
    assign mux_in_cos106 = 16'b0010001000100100;
    assign mux_in_sin106 = 16'b0111101101011101;
    assign mux_in_cos107 = 16'b0010000010011111;
    assign mux_in_sin107 = 16'b0111101111000110;
    assign mux_in_cos108 = 16'b0001111100011010;
    assign mux_in_sin108 = 16'b0111110000101010;
    assign mux_in_cos109 = 16'b0001110110010011;
    assign mux_in_sin109 = 16'b0111110010001001;
    assign mux_in_cos110 = 16'b0001110000001100;
    assign mux_in_sin110 = 16'b0111110011100100;
    assign mux_in_cos111 = 16'b0001101010000011;
    assign mux_in_sin111 = 16'b0111110100111010;
    assign mux_in_cos112 = 16'b0001100011111001;
    assign mux_in_sin112 = 16'b0111110110001010;
    assign mux_in_cos113 = 16'b0001011101101110;
    assign mux_in_sin113 = 16'b0111110111010110;
    assign mux_in_cos114 = 16'b0001010111100010;
    assign mux_in_sin114 = 16'b0111111000011110;
    assign mux_in_cos115 = 16'b0001010001010101;
    assign mux_in_sin115 = 16'b0111111001100000;
    assign mux_in_cos116 = 16'b0001001011001000;
    assign mux_in_sin116 = 16'b0111111010011101;
    assign mux_in_cos117 = 16'b0001000100111010;
    assign mux_in_sin117 = 16'b0111111011010110;
    assign mux_in_cos118 = 16'b0000111110101011;
    assign mux_in_sin118 = 16'b0111111100001010;
    assign mux_in_cos119 = 16'b0000111000011100;
    assign mux_in_sin119 = 16'b0111111100111000;
    assign mux_in_cos120 = 16'b0000110010001100;
    assign mux_in_sin120 = 16'b0111111101100010;
    assign mux_in_cos121 = 16'b0000101011111011;
    assign mux_in_sin121 = 16'b0111111110000111;
    assign mux_in_cos122 = 16'b0000100101101011;
    assign mux_in_sin122 = 16'b0111111110100111;
    assign mux_in_cos123 = 16'b0000011111011001;
    assign mux_in_sin123 = 16'b0111111111000010;
    assign mux_in_cos124 = 16'b0000011001001000;
    assign mux_in_sin124 = 16'b0111111111011001;
    assign mux_in_cos125 = 16'b0000010010110110;
    assign mux_in_sin125 = 16'b0111111111101010;
    assign mux_in_cos126 = 16'b0000001100100100;
    assign mux_in_sin126 = 16'b0111111111110110;
    assign mux_in_cos127 = 16'b0000000110010010;
    assign mux_in_sin127 = 16'b0111111111111110;
    assign mux_in_cos128 = 16'b0000000000000000;
    assign mux_in_sin128 = 16'b1000000000000000;

    // Sine LUTs

    always @ (*)
    begin
        case(x_in1)
        8'b00000000 : sin1 = mux_in_sin0;
        8'b00000001 : sin1 = mux_in_sin1;
        8'b00000010 : sin1 = mux_in_sin2;
        8'b00000011 : sin1 = mux_in_sin3;
        8'b00000100 : sin1 = mux_in_sin4;
        8'b00000101 : sin1 = mux_in_sin5;
        8'b00000110 : sin1 = mux_in_sin6;
        8'b00000111 : sin1 = mux_in_sin7;
        8'b00001000 : sin1 = mux_in_sin8;
        8'b00001001 : sin1 = mux_in_sin9;
        8'b00001010 : sin1 = mux_in_sin10;
        8'b00001011 : sin1 = mux_in_sin11;
        8'b00001100 : sin1 = mux_in_sin12;
        8'b00001101 : sin1 = mux_in_sin13;
        8'b00001110 : sin1 = mux_in_sin14;
        8'b00001111 : sin1 = mux_in_sin15;
        8'b00010000 : sin1 = mux_in_sin16;
        8'b00010001 : sin1 = mux_in_sin17;
        8'b00010010 : sin1 = mux_in_sin18;
        8'b00010011 : sin1 = mux_in_sin19;
        8'b00010100 : sin1 = mux_in_sin20;
        8'b00010101 : sin1 = mux_in_sin21;
        8'b00010110 : sin1 = mux_in_sin22;
        8'b00010111 : sin1 = mux_in_sin23;
        8'b00011000 : sin1 = mux_in_sin24;
        8'b00011001 : sin1 = mux_in_sin25;
        8'b00011010 : sin1 = mux_in_sin26;
        8'b00011011 : sin1 = mux_in_sin27;
        8'b00011100 : sin1 = mux_in_sin28;
        8'b00011101 : sin1 = mux_in_sin29;
        8'b00011110 : sin1 = mux_in_sin30;
        8'b00011111 : sin1 = mux_in_sin31;
        8'b00100000 : sin1 = mux_in_sin32;
        8'b00100001 : sin1 = mux_in_sin33;
        8'b00100010 : sin1 = mux_in_sin34;
        8'b00100011 : sin1 = mux_in_sin35;
        8'b00100100 : sin1 = mux_in_sin36;
        8'b00100101 : sin1 = mux_in_sin37;
        8'b00100110 : sin1 = mux_in_sin38;
        8'b00100111 : sin1 = mux_in_sin39;
        8'b00101000 : sin1 = mux_in_sin40;
        8'b00101001 : sin1 = mux_in_sin41;
        8'b00101010 : sin1 = mux_in_sin42;
        8'b00101011 : sin1 = mux_in_sin43;
        8'b00101100 : sin1 = mux_in_sin44;
        8'b00101101 : sin1 = mux_in_sin45;
        8'b00101110 : sin1 = mux_in_sin46;
        8'b00101111 : sin1 = mux_in_sin47;
        8'b00110000 : sin1 = mux_in_sin48;
        8'b00110001 : sin1 = mux_in_sin49;
        8'b00110010 : sin1 = mux_in_sin50;
        8'b00110011 : sin1 = mux_in_sin51;
        8'b00110100 : sin1 = mux_in_sin52;
        8'b00110101 : sin1 = mux_in_sin53;
        8'b00110110 : sin1 = mux_in_sin54;
        8'b00110111 : sin1 = mux_in_sin55;
        8'b00111000 : sin1 = mux_in_sin56;
        8'b00111001 : sin1 = mux_in_sin57;
        8'b00111010 : sin1 = mux_in_sin58;
        8'b00111011 : sin1 = mux_in_sin59;
        8'b00111100 : sin1 = mux_in_sin60;
        8'b00111101 : sin1 = mux_in_sin61;
        8'b00111110 : sin1 = mux_in_sin62;
        8'b00111111 : sin1 = mux_in_sin63;
        8'b01000000 : sin1 = mux_in_sin64;
        8'b01000001 : sin1 = mux_in_sin65;
        8'b01000010 : sin1 = mux_in_sin66;
        8'b01000011 : sin1 = mux_in_sin67;
        8'b01000100 : sin1 = mux_in_sin68;
        8'b01000101 : sin1 = mux_in_sin69;
        8'b01000110 : sin1 = mux_in_sin70;
        8'b01000111 : sin1 = mux_in_sin71;
        8'b01001000 : sin1 = mux_in_sin72;
        8'b01001001 : sin1 = mux_in_sin73;
        8'b01001010 : sin1 = mux_in_sin74;
        8'b01001011 : sin1 = mux_in_sin75;
        8'b01001100 : sin1 = mux_in_sin76;
        8'b01001101 : sin1 = mux_in_sin77;
        8'b01001110 : sin1 = mux_in_sin78;
        8'b01001111 : sin1 = mux_in_sin79;
        8'b01010000 : sin1 = mux_in_sin80;
        8'b01010001 : sin1 = mux_in_sin81;
        8'b01010010 : sin1 = mux_in_sin82;
        8'b01010011 : sin1 = mux_in_sin83;
        8'b01010100 : sin1 = mux_in_sin84;
        8'b01010101 : sin1 = mux_in_sin85;
        8'b01010110 : sin1 = mux_in_sin86;
        8'b01010111 : sin1 = mux_in_sin87;
        8'b01011000 : sin1 = mux_in_sin88;
        8'b01011001 : sin1 = mux_in_sin89;
        8'b01011010 : sin1 = mux_in_sin90;
        8'b01011011 : sin1 = mux_in_sin91;
        8'b01011100 : sin1 = mux_in_sin92;
        8'b01011101 : sin1 = mux_in_sin93;
        8'b01011110 : sin1 = mux_in_sin94;
        8'b01011111 : sin1 = mux_in_sin95;
        8'b01100000 : sin1 = mux_in_sin96;
        8'b01100001 : sin1 = mux_in_sin97;
        8'b01100010 : sin1 = mux_in_sin98;
        8'b01100011 : sin1 = mux_in_sin99;
        8'b01100100 : sin1 = mux_in_sin100;
        8'b01100101 : sin1 = mux_in_sin101;
        8'b01100110 : sin1 = mux_in_sin102;
        8'b01100111 : sin1 = mux_in_sin103;
        8'b01101000 : sin1 = mux_in_sin104;
        8'b01101001 : sin1 = mux_in_sin105;
        8'b01101010 : sin1 = mux_in_sin106;
        8'b01101011 : sin1 = mux_in_sin107;
        8'b01101100 : sin1 = mux_in_sin108;
        8'b01101101 : sin1 = mux_in_sin109;
        8'b01101110 : sin1 = mux_in_sin110;
        8'b01101111 : sin1 = mux_in_sin111;
        8'b01110000 : sin1 = mux_in_sin112;
        8'b01110001 : sin1 = mux_in_sin113;
        8'b01110010 : sin1 = mux_in_sin114;
        8'b01110011 : sin1 = mux_in_sin115;
        8'b01110100 : sin1 = mux_in_sin116;
        8'b01110101 : sin1 = mux_in_sin117;
        8'b01110110 : sin1 = mux_in_sin118;
        8'b01110111 : sin1 = mux_in_sin119;
        8'b01111000 : sin1 = mux_in_sin120;
        8'b01111001 : sin1 = mux_in_sin121;
        8'b01111010 : sin1 = mux_in_sin122;
        8'b01111011 : sin1 = mux_in_sin123;
        8'b01111100 : sin1 = mux_in_sin124;
        8'b01111101 : sin1 = mux_in_sin125;
        8'b01111110 : sin1 = mux_in_sin126;
        8'b01111111 : sin1 = mux_in_sin127;
        8'b10000000 : sin1 = mux_in_sin128;
        default: sin1 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in2)
        8'b00000000 : sin2 = mux_in_sin0;
        8'b00000001 : sin2 = mux_in_sin1;
        8'b00000010 : sin2 = mux_in_sin2;
        8'b00000011 : sin2 = mux_in_sin3;
        8'b00000100 : sin2 = mux_in_sin4;
        8'b00000101 : sin2 = mux_in_sin5;
        8'b00000110 : sin2 = mux_in_sin6;
        8'b00000111 : sin2 = mux_in_sin7;
        8'b00001000 : sin2 = mux_in_sin8;
        8'b00001001 : sin2 = mux_in_sin9;
        8'b00001010 : sin2 = mux_in_sin10;
        8'b00001011 : sin2 = mux_in_sin11;
        8'b00001100 : sin2 = mux_in_sin12;
        8'b00001101 : sin2 = mux_in_sin13;
        8'b00001110 : sin2 = mux_in_sin14;
        8'b00001111 : sin2 = mux_in_sin15;
        8'b00010000 : sin2 = mux_in_sin16;
        8'b00010001 : sin2 = mux_in_sin17;
        8'b00010010 : sin2 = mux_in_sin18;
        8'b00010011 : sin2 = mux_in_sin19;
        8'b00010100 : sin2 = mux_in_sin20;
        8'b00010101 : sin2 = mux_in_sin21;
        8'b00010110 : sin2 = mux_in_sin22;
        8'b00010111 : sin2 = mux_in_sin23;
        8'b00011000 : sin2 = mux_in_sin24;
        8'b00011001 : sin2 = mux_in_sin25;
        8'b00011010 : sin2 = mux_in_sin26;
        8'b00011011 : sin2 = mux_in_sin27;
        8'b00011100 : sin2 = mux_in_sin28;
        8'b00011101 : sin2 = mux_in_sin29;
        8'b00011110 : sin2 = mux_in_sin30;
        8'b00011111 : sin2 = mux_in_sin31;
        8'b00100000 : sin2 = mux_in_sin32;
        8'b00100001 : sin2 = mux_in_sin33;
        8'b00100010 : sin2 = mux_in_sin34;
        8'b00100011 : sin2 = mux_in_sin35;
        8'b00100100 : sin2 = mux_in_sin36;
        8'b00100101 : sin2 = mux_in_sin37;
        8'b00100110 : sin2 = mux_in_sin38;
        8'b00100111 : sin2 = mux_in_sin39;
        8'b00101000 : sin2 = mux_in_sin40;
        8'b00101001 : sin2 = mux_in_sin41;
        8'b00101010 : sin2 = mux_in_sin42;
        8'b00101011 : sin2 = mux_in_sin43;
        8'b00101100 : sin2 = mux_in_sin44;
        8'b00101101 : sin2 = mux_in_sin45;
        8'b00101110 : sin2 = mux_in_sin46;
        8'b00101111 : sin2 = mux_in_sin47;
        8'b00110000 : sin2 = mux_in_sin48;
        8'b00110001 : sin2 = mux_in_sin49;
        8'b00110010 : sin2 = mux_in_sin50;
        8'b00110011 : sin2 = mux_in_sin51;
        8'b00110100 : sin2 = mux_in_sin52;
        8'b00110101 : sin2 = mux_in_sin53;
        8'b00110110 : sin2 = mux_in_sin54;
        8'b00110111 : sin2 = mux_in_sin55;
        8'b00111000 : sin2 = mux_in_sin56;
        8'b00111001 : sin2 = mux_in_sin57;
        8'b00111010 : sin2 = mux_in_sin58;
        8'b00111011 : sin2 = mux_in_sin59;
        8'b00111100 : sin2 = mux_in_sin60;
        8'b00111101 : sin2 = mux_in_sin61;
        8'b00111110 : sin2 = mux_in_sin62;
        8'b00111111 : sin2 = mux_in_sin63;
        8'b01000000 : sin2 = mux_in_sin64;
        8'b01000001 : sin2 = mux_in_sin65;
        8'b01000010 : sin2 = mux_in_sin66;
        8'b01000011 : sin2 = mux_in_sin67;
        8'b01000100 : sin2 = mux_in_sin68;
        8'b01000101 : sin2 = mux_in_sin69;
        8'b01000110 : sin2 = mux_in_sin70;
        8'b01000111 : sin2 = mux_in_sin71;
        8'b01001000 : sin2 = mux_in_sin72;
        8'b01001001 : sin2 = mux_in_sin73;
        8'b01001010 : sin2 = mux_in_sin74;
        8'b01001011 : sin2 = mux_in_sin75;
        8'b01001100 : sin2 = mux_in_sin76;
        8'b01001101 : sin2 = mux_in_sin77;
        8'b01001110 : sin2 = mux_in_sin78;
        8'b01001111 : sin2 = mux_in_sin79;
        8'b01010000 : sin2 = mux_in_sin80;
        8'b01010001 : sin2 = mux_in_sin81;
        8'b01010010 : sin2 = mux_in_sin82;
        8'b01010011 : sin2 = mux_in_sin83;
        8'b01010100 : sin2 = mux_in_sin84;
        8'b01010101 : sin2 = mux_in_sin85;
        8'b01010110 : sin2 = mux_in_sin86;
        8'b01010111 : sin2 = mux_in_sin87;
        8'b01011000 : sin2 = mux_in_sin88;
        8'b01011001 : sin2 = mux_in_sin89;
        8'b01011010 : sin2 = mux_in_sin90;
        8'b01011011 : sin2 = mux_in_sin91;
        8'b01011100 : sin2 = mux_in_sin92;
        8'b01011101 : sin2 = mux_in_sin93;
        8'b01011110 : sin2 = mux_in_sin94;
        8'b01011111 : sin2 = mux_in_sin95;
        8'b01100000 : sin2 = mux_in_sin96;
        8'b01100001 : sin2 = mux_in_sin97;
        8'b01100010 : sin2 = mux_in_sin98;
        8'b01100011 : sin2 = mux_in_sin99;
        8'b01100100 : sin2 = mux_in_sin100;
        8'b01100101 : sin2 = mux_in_sin101;
        8'b01100110 : sin2 = mux_in_sin102;
        8'b01100111 : sin2 = mux_in_sin103;
        8'b01101000 : sin2 = mux_in_sin104;
        8'b01101001 : sin2 = mux_in_sin105;
        8'b01101010 : sin2 = mux_in_sin106;
        8'b01101011 : sin2 = mux_in_sin107;
        8'b01101100 : sin2 = mux_in_sin108;
        8'b01101101 : sin2 = mux_in_sin109;
        8'b01101110 : sin2 = mux_in_sin110;
        8'b01101111 : sin2 = mux_in_sin111;
        8'b01110000 : sin2 = mux_in_sin112;
        8'b01110001 : sin2 = mux_in_sin113;
        8'b01110010 : sin2 = mux_in_sin114;
        8'b01110011 : sin2 = mux_in_sin115;
        8'b01110100 : sin2 = mux_in_sin116;
        8'b01110101 : sin2 = mux_in_sin117;
        8'b01110110 : sin2 = mux_in_sin118;
        8'b01110111 : sin2 = mux_in_sin119;
        8'b01111000 : sin2 = mux_in_sin120;
        8'b01111001 : sin2 = mux_in_sin121;
        8'b01111010 : sin2 = mux_in_sin122;
        8'b01111011 : sin2 = mux_in_sin123;
        8'b01111100 : sin2 = mux_in_sin124;
        8'b01111101 : sin2 = mux_in_sin125;
        8'b01111110 : sin2 = mux_in_sin126;
        8'b01111111 : sin2 = mux_in_sin127;
        8'b10000000 : sin2 = mux_in_sin128;
        default: sin2 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in3)
        8'b00000000 : sin3 = mux_in_sin0;
        8'b00000001 : sin3 = mux_in_sin1;
        8'b00000010 : sin3 = mux_in_sin2;
        8'b00000011 : sin3 = mux_in_sin3;
        8'b00000100 : sin3 = mux_in_sin4;
        8'b00000101 : sin3 = mux_in_sin5;
        8'b00000110 : sin3 = mux_in_sin6;
        8'b00000111 : sin3 = mux_in_sin7;
        8'b00001000 : sin3 = mux_in_sin8;
        8'b00001001 : sin3 = mux_in_sin9;
        8'b00001010 : sin3 = mux_in_sin10;
        8'b00001011 : sin3 = mux_in_sin11;
        8'b00001100 : sin3 = mux_in_sin12;
        8'b00001101 : sin3 = mux_in_sin13;
        8'b00001110 : sin3 = mux_in_sin14;
        8'b00001111 : sin3 = mux_in_sin15;
        8'b00010000 : sin3 = mux_in_sin16;
        8'b00010001 : sin3 = mux_in_sin17;
        8'b00010010 : sin3 = mux_in_sin18;
        8'b00010011 : sin3 = mux_in_sin19;
        8'b00010100 : sin3 = mux_in_sin20;
        8'b00010101 : sin3 = mux_in_sin21;
        8'b00010110 : sin3 = mux_in_sin22;
        8'b00010111 : sin3 = mux_in_sin23;
        8'b00011000 : sin3 = mux_in_sin24;
        8'b00011001 : sin3 = mux_in_sin25;
        8'b00011010 : sin3 = mux_in_sin26;
        8'b00011011 : sin3 = mux_in_sin27;
        8'b00011100 : sin3 = mux_in_sin28;
        8'b00011101 : sin3 = mux_in_sin29;
        8'b00011110 : sin3 = mux_in_sin30;
        8'b00011111 : sin3 = mux_in_sin31;
        8'b00100000 : sin3 = mux_in_sin32;
        8'b00100001 : sin3 = mux_in_sin33;
        8'b00100010 : sin3 = mux_in_sin34;
        8'b00100011 : sin3 = mux_in_sin35;
        8'b00100100 : sin3 = mux_in_sin36;
        8'b00100101 : sin3 = mux_in_sin37;
        8'b00100110 : sin3 = mux_in_sin38;
        8'b00100111 : sin3 = mux_in_sin39;
        8'b00101000 : sin3 = mux_in_sin40;
        8'b00101001 : sin3 = mux_in_sin41;
        8'b00101010 : sin3 = mux_in_sin42;
        8'b00101011 : sin3 = mux_in_sin43;
        8'b00101100 : sin3 = mux_in_sin44;
        8'b00101101 : sin3 = mux_in_sin45;
        8'b00101110 : sin3 = mux_in_sin46;
        8'b00101111 : sin3 = mux_in_sin47;
        8'b00110000 : sin3 = mux_in_sin48;
        8'b00110001 : sin3 = mux_in_sin49;
        8'b00110010 : sin3 = mux_in_sin50;
        8'b00110011 : sin3 = mux_in_sin51;
        8'b00110100 : sin3 = mux_in_sin52;
        8'b00110101 : sin3 = mux_in_sin53;
        8'b00110110 : sin3 = mux_in_sin54;
        8'b00110111 : sin3 = mux_in_sin55;
        8'b00111000 : sin3 = mux_in_sin56;
        8'b00111001 : sin3 = mux_in_sin57;
        8'b00111010 : sin3 = mux_in_sin58;
        8'b00111011 : sin3 = mux_in_sin59;
        8'b00111100 : sin3 = mux_in_sin60;
        8'b00111101 : sin3 = mux_in_sin61;
        8'b00111110 : sin3 = mux_in_sin62;
        8'b00111111 : sin3 = mux_in_sin63;
        8'b01000000 : sin3 = mux_in_sin64;
        8'b01000001 : sin3 = mux_in_sin65;
        8'b01000010 : sin3 = mux_in_sin66;
        8'b01000011 : sin3 = mux_in_sin67;
        8'b01000100 : sin3 = mux_in_sin68;
        8'b01000101 : sin3 = mux_in_sin69;
        8'b01000110 : sin3 = mux_in_sin70;
        8'b01000111 : sin3 = mux_in_sin71;
        8'b01001000 : sin3 = mux_in_sin72;
        8'b01001001 : sin3 = mux_in_sin73;
        8'b01001010 : sin3 = mux_in_sin74;
        8'b01001011 : sin3 = mux_in_sin75;
        8'b01001100 : sin3 = mux_in_sin76;
        8'b01001101 : sin3 = mux_in_sin77;
        8'b01001110 : sin3 = mux_in_sin78;
        8'b01001111 : sin3 = mux_in_sin79;
        8'b01010000 : sin3 = mux_in_sin80;
        8'b01010001 : sin3 = mux_in_sin81;
        8'b01010010 : sin3 = mux_in_sin82;
        8'b01010011 : sin3 = mux_in_sin83;
        8'b01010100 : sin3 = mux_in_sin84;
        8'b01010101 : sin3 = mux_in_sin85;
        8'b01010110 : sin3 = mux_in_sin86;
        8'b01010111 : sin3 = mux_in_sin87;
        8'b01011000 : sin3 = mux_in_sin88;
        8'b01011001 : sin3 = mux_in_sin89;
        8'b01011010 : sin3 = mux_in_sin90;
        8'b01011011 : sin3 = mux_in_sin91;
        8'b01011100 : sin3 = mux_in_sin92;
        8'b01011101 : sin3 = mux_in_sin93;
        8'b01011110 : sin3 = mux_in_sin94;
        8'b01011111 : sin3 = mux_in_sin95;
        8'b01100000 : sin3 = mux_in_sin96;
        8'b01100001 : sin3 = mux_in_sin97;
        8'b01100010 : sin3 = mux_in_sin98;
        8'b01100011 : sin3 = mux_in_sin99;
        8'b01100100 : sin3 = mux_in_sin100;
        8'b01100101 : sin3 = mux_in_sin101;
        8'b01100110 : sin3 = mux_in_sin102;
        8'b01100111 : sin3 = mux_in_sin103;
        8'b01101000 : sin3 = mux_in_sin104;
        8'b01101001 : sin3 = mux_in_sin105;
        8'b01101010 : sin3 = mux_in_sin106;
        8'b01101011 : sin3 = mux_in_sin107;
        8'b01101100 : sin3 = mux_in_sin108;
        8'b01101101 : sin3 = mux_in_sin109;
        8'b01101110 : sin3 = mux_in_sin110;
        8'b01101111 : sin3 = mux_in_sin111;
        8'b01110000 : sin3 = mux_in_sin112;
        8'b01110001 : sin3 = mux_in_sin113;
        8'b01110010 : sin3 = mux_in_sin114;
        8'b01110011 : sin3 = mux_in_sin115;
        8'b01110100 : sin3 = mux_in_sin116;
        8'b01110101 : sin3 = mux_in_sin117;
        8'b01110110 : sin3 = mux_in_sin118;
        8'b01110111 : sin3 = mux_in_sin119;
        8'b01111000 : sin3 = mux_in_sin120;
        8'b01111001 : sin3 = mux_in_sin121;
        8'b01111010 : sin3 = mux_in_sin122;
        8'b01111011 : sin3 = mux_in_sin123;
        8'b01111100 : sin3 = mux_in_sin124;
        8'b01111101 : sin3 = mux_in_sin125;
        8'b01111110 : sin3 = mux_in_sin126;
        8'b01111111 : sin3 = mux_in_sin127;
        8'b10000000 : sin3 = mux_in_sin128;
        default: sin3 = 15'bx;
        endcase
    end

    //Cos LUTs
    always @ (*)
    begin
        case(x_in1)
        8'b00000000 : cos1 = mux_in_cos0;
        8'b00000001 : cos1 = mux_in_cos1;
        8'b00000010 : cos1 = mux_in_cos2;
        8'b00000011 : cos1 = mux_in_cos3;
        8'b00000100 : cos1 = mux_in_cos4;
        8'b00000101 : cos1 = mux_in_cos5;
        8'b00000110 : cos1 = mux_in_cos6;
        8'b00000111 : cos1 = mux_in_cos7;
        8'b00001000 : cos1 = mux_in_cos8;
        8'b00001001 : cos1 = mux_in_cos9;
        8'b00001010 : cos1 = mux_in_cos10;
        8'b00001011 : cos1 = mux_in_cos11;
        8'b00001100 : cos1 = mux_in_cos12;
        8'b00001101 : cos1 = mux_in_cos13;
        8'b00001110 : cos1 = mux_in_cos14;
        8'b00001111 : cos1 = mux_in_cos15;
        8'b00010000 : cos1 = mux_in_cos16;
        8'b00010001 : cos1 = mux_in_cos17;
        8'b00010010 : cos1 = mux_in_cos18;
        8'b00010011 : cos1 = mux_in_cos19;
        8'b00010100 : cos1 = mux_in_cos20;
        8'b00010101 : cos1 = mux_in_cos21;
        8'b00010110 : cos1 = mux_in_cos22;
        8'b00010111 : cos1 = mux_in_cos23;
        8'b00011000 : cos1 = mux_in_cos24;
        8'b00011001 : cos1 = mux_in_cos25;
        8'b00011010 : cos1 = mux_in_cos26;
        8'b00011011 : cos1 = mux_in_cos27;
        8'b00011100 : cos1 = mux_in_cos28;
        8'b00011101 : cos1 = mux_in_cos29;
        8'b00011110 : cos1 = mux_in_cos30;
        8'b00011111 : cos1 = mux_in_cos31;
        8'b00100000 : cos1 = mux_in_cos32;
        8'b00100001 : cos1 = mux_in_cos33;
        8'b00100010 : cos1 = mux_in_cos34;
        8'b00100011 : cos1 = mux_in_cos35;
        8'b00100100 : cos1 = mux_in_cos36;
        8'b00100101 : cos1 = mux_in_cos37;
        8'b00100110 : cos1 = mux_in_cos38;
        8'b00100111 : cos1 = mux_in_cos39;
        8'b00101000 : cos1 = mux_in_cos40;
        8'b00101001 : cos1 = mux_in_cos41;
        8'b00101010 : cos1 = mux_in_cos42;
        8'b00101011 : cos1 = mux_in_cos43;
        8'b00101100 : cos1 = mux_in_cos44;
        8'b00101101 : cos1 = mux_in_cos45;
        8'b00101110 : cos1 = mux_in_cos46;
        8'b00101111 : cos1 = mux_in_cos47;
        8'b00110000 : cos1 = mux_in_cos48;
        8'b00110001 : cos1 = mux_in_cos49;
        8'b00110010 : cos1 = mux_in_cos50;
        8'b00110011 : cos1 = mux_in_cos51;
        8'b00110100 : cos1 = mux_in_cos52;
        8'b00110101 : cos1 = mux_in_cos53;
        8'b00110110 : cos1 = mux_in_cos54;
        8'b00110111 : cos1 = mux_in_cos55;
        8'b00111000 : cos1 = mux_in_cos56;
        8'b00111001 : cos1 = mux_in_cos57;
        8'b00111010 : cos1 = mux_in_cos58;
        8'b00111011 : cos1 = mux_in_cos59;
        8'b00111100 : cos1 = mux_in_cos60;
        8'b00111101 : cos1 = mux_in_cos61;
        8'b00111110 : cos1 = mux_in_cos62;
        8'b00111111 : cos1 = mux_in_cos63;
        8'b01000000 : cos1 = mux_in_cos64;
        8'b01000001 : cos1 = mux_in_cos65;
        8'b01000010 : cos1 = mux_in_cos66;
        8'b01000011 : cos1 = mux_in_cos67;
        8'b01000100 : cos1 = mux_in_cos68;
        8'b01000101 : cos1 = mux_in_cos69;
        8'b01000110 : cos1 = mux_in_cos70;
        8'b01000111 : cos1 = mux_in_cos71;
        8'b01001000 : cos1 = mux_in_cos72;
        8'b01001001 : cos1 = mux_in_cos73;
        8'b01001010 : cos1 = mux_in_cos74;
        8'b01001011 : cos1 = mux_in_cos75;
        8'b01001100 : cos1 = mux_in_cos76;
        8'b01001101 : cos1 = mux_in_cos77;
        8'b01001110 : cos1 = mux_in_cos78;
        8'b01001111 : cos1 = mux_in_cos79;
        8'b01010000 : cos1 = mux_in_cos80;
        8'b01010001 : cos1 = mux_in_cos81;
        8'b01010010 : cos1 = mux_in_cos82;
        8'b01010011 : cos1 = mux_in_cos83;
        8'b01010100 : cos1 = mux_in_cos84;
        8'b01010101 : cos1 = mux_in_cos85;
        8'b01010110 : cos1 = mux_in_cos86;
        8'b01010111 : cos1 = mux_in_cos87;
        8'b01011000 : cos1 = mux_in_cos88;
        8'b01011001 : cos1 = mux_in_cos89;
        8'b01011010 : cos1 = mux_in_cos90;
        8'b01011011 : cos1 = mux_in_cos91;
        8'b01011100 : cos1 = mux_in_cos92;
        8'b01011101 : cos1 = mux_in_cos93;
        8'b01011110 : cos1 = mux_in_cos94;
        8'b01011111 : cos1 = mux_in_cos95;
        8'b01100000 : cos1 = mux_in_cos96;
        8'b01100001 : cos1 = mux_in_cos97;
        8'b01100010 : cos1 = mux_in_cos98;
        8'b01100011 : cos1 = mux_in_cos99;
        8'b01100100 : cos1 = mux_in_cos100;
        8'b01100101 : cos1 = mux_in_cos101;
        8'b01100110 : cos1 = mux_in_cos102;
        8'b01100111 : cos1 = mux_in_cos103;
        8'b01101000 : cos1 = mux_in_cos104;
        8'b01101001 : cos1 = mux_in_cos105;
        8'b01101010 : cos1 = mux_in_cos106;
        8'b01101011 : cos1 = mux_in_cos107;
        8'b01101100 : cos1 = mux_in_cos108;
        8'b01101101 : cos1 = mux_in_cos109;
        8'b01101110 : cos1 = mux_in_cos110;
        8'b01101111 : cos1 = mux_in_cos111;
        8'b01110000 : cos1 = mux_in_cos112;
        8'b01110001 : cos1 = mux_in_cos113;
        8'b01110010 : cos1 = mux_in_cos114;
        8'b01110011 : cos1 = mux_in_cos115;
        8'b01110100 : cos1 = mux_in_cos116;
        8'b01110101 : cos1 = mux_in_cos117;
        8'b01110110 : cos1 = mux_in_cos118;
        8'b01110111 : cos1 = mux_in_cos119;
        8'b01111000 : cos1 = mux_in_cos120;
        8'b01111001 : cos1 = mux_in_cos121;
        8'b01111010 : cos1 = mux_in_cos122;
        8'b01111011 : cos1 = mux_in_cos123;
        8'b01111100 : cos1 = mux_in_cos124;
        8'b01111101 : cos1 = mux_in_cos125;
        8'b01111110 : cos1 = mux_in_cos126;
        8'b01111111 : cos1 = mux_in_cos127;
        8'b10000000 : cos1 = mux_in_cos128;
        default: cos1 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in2)
        8'b00000000 : cos2 = mux_in_cos0;
        8'b00000001 : cos2 = mux_in_cos1;
        8'b00000010 : cos2 = mux_in_cos2;
        8'b00000011 : cos2 = mux_in_cos3;
        8'b00000100 : cos2 = mux_in_cos4;
        8'b00000101 : cos2 = mux_in_cos5;
        8'b00000110 : cos2 = mux_in_cos6;
        8'b00000111 : cos2 = mux_in_cos7;
        8'b00001000 : cos2 = mux_in_cos8;
        8'b00001001 : cos2 = mux_in_cos9;
        8'b00001010 : cos2 = mux_in_cos10;
        8'b00001011 : cos2 = mux_in_cos11;
        8'b00001100 : cos2 = mux_in_cos12;
        8'b00001101 : cos2 = mux_in_cos13;
        8'b00001110 : cos2 = mux_in_cos14;
        8'b00001111 : cos2 = mux_in_cos15;
        8'b00010000 : cos2 = mux_in_cos16;
        8'b00010001 : cos2 = mux_in_cos17;
        8'b00010010 : cos2 = mux_in_cos18;
        8'b00010011 : cos2 = mux_in_cos19;
        8'b00010100 : cos2 = mux_in_cos20;
        8'b00010101 : cos2 = mux_in_cos21;
        8'b00010110 : cos2 = mux_in_cos22;
        8'b00010111 : cos2 = mux_in_cos23;
        8'b00011000 : cos2 = mux_in_cos24;
        8'b00011001 : cos2 = mux_in_cos25;
        8'b00011010 : cos2 = mux_in_cos26;
        8'b00011011 : cos2 = mux_in_cos27;
        8'b00011100 : cos2 = mux_in_cos28;
        8'b00011101 : cos2 = mux_in_cos29;
        8'b00011110 : cos2 = mux_in_cos30;
        8'b00011111 : cos2 = mux_in_cos31;
        8'b00100000 : cos2 = mux_in_cos32;
        8'b00100001 : cos2 = mux_in_cos33;
        8'b00100010 : cos2 = mux_in_cos34;
        8'b00100011 : cos2 = mux_in_cos35;
        8'b00100100 : cos2 = mux_in_cos36;
        8'b00100101 : cos2 = mux_in_cos37;
        8'b00100110 : cos2 = mux_in_cos38;
        8'b00100111 : cos2 = mux_in_cos39;
        8'b00101000 : cos2 = mux_in_cos40;
        8'b00101001 : cos2 = mux_in_cos41;
        8'b00101010 : cos2 = mux_in_cos42;
        8'b00101011 : cos2 = mux_in_cos43;
        8'b00101100 : cos2 = mux_in_cos44;
        8'b00101101 : cos2 = mux_in_cos45;
        8'b00101110 : cos2 = mux_in_cos46;
        8'b00101111 : cos2 = mux_in_cos47;
        8'b00110000 : cos2 = mux_in_cos48;
        8'b00110001 : cos2 = mux_in_cos49;
        8'b00110010 : cos2 = mux_in_cos50;
        8'b00110011 : cos2 = mux_in_cos51;
        8'b00110100 : cos2 = mux_in_cos52;
        8'b00110101 : cos2 = mux_in_cos53;
        8'b00110110 : cos2 = mux_in_cos54;
        8'b00110111 : cos2 = mux_in_cos55;
        8'b00111000 : cos2 = mux_in_cos56;
        8'b00111001 : cos2 = mux_in_cos57;
        8'b00111010 : cos2 = mux_in_cos58;
        8'b00111011 : cos2 = mux_in_cos59;
        8'b00111100 : cos2 = mux_in_cos60;
        8'b00111101 : cos2 = mux_in_cos61;
        8'b00111110 : cos2 = mux_in_cos62;
        8'b00111111 : cos2 = mux_in_cos63;
        8'b01000000 : cos2 = mux_in_cos64;
        8'b01000001 : cos2 = mux_in_cos65;
        8'b01000010 : cos2 = mux_in_cos66;
        8'b01000011 : cos2 = mux_in_cos67;
        8'b01000100 : cos2 = mux_in_cos68;
        8'b01000101 : cos2 = mux_in_cos69;
        8'b01000110 : cos2 = mux_in_cos70;
        8'b01000111 : cos2 = mux_in_cos71;
        8'b01001000 : cos2 = mux_in_cos72;
        8'b01001001 : cos2 = mux_in_cos73;
        8'b01001010 : cos2 = mux_in_cos74;
        8'b01001011 : cos2 = mux_in_cos75;
        8'b01001100 : cos2 = mux_in_cos76;
        8'b01001101 : cos2 = mux_in_cos77;
        8'b01001110 : cos2 = mux_in_cos78;
        8'b01001111 : cos2 = mux_in_cos79;
        8'b01010000 : cos2 = mux_in_cos80;
        8'b01010001 : cos2 = mux_in_cos81;
        8'b01010010 : cos2 = mux_in_cos82;
        8'b01010011 : cos2 = mux_in_cos83;
        8'b01010100 : cos2 = mux_in_cos84;
        8'b01010101 : cos2 = mux_in_cos85;
        8'b01010110 : cos2 = mux_in_cos86;
        8'b01010111 : cos2 = mux_in_cos87;
        8'b01011000 : cos2 = mux_in_cos88;
        8'b01011001 : cos2 = mux_in_cos89;
        8'b01011010 : cos2 = mux_in_cos90;
        8'b01011011 : cos2 = mux_in_cos91;
        8'b01011100 : cos2 = mux_in_cos92;
        8'b01011101 : cos2 = mux_in_cos93;
        8'b01011110 : cos2 = mux_in_cos94;
        8'b01011111 : cos2 = mux_in_cos95;
        8'b01100000 : cos2 = mux_in_cos96;
        8'b01100001 : cos2 = mux_in_cos97;
        8'b01100010 : cos2 = mux_in_cos98;
        8'b01100011 : cos2 = mux_in_cos99;
        8'b01100100 : cos2 = mux_in_cos100;
        8'b01100101 : cos2 = mux_in_cos101;
        8'b01100110 : cos2 = mux_in_cos102;
        8'b01100111 : cos2 = mux_in_cos103;
        8'b01101000 : cos2 = mux_in_cos104;
        8'b01101001 : cos2 = mux_in_cos105;
        8'b01101010 : cos2 = mux_in_cos106;
        8'b01101011 : cos2 = mux_in_cos107;
        8'b01101100 : cos2 = mux_in_cos108;
        8'b01101101 : cos2 = mux_in_cos109;
        8'b01101110 : cos2 = mux_in_cos110;
        8'b01101111 : cos2 = mux_in_cos111;
        8'b01110000 : cos2 = mux_in_cos112;
        8'b01110001 : cos2 = mux_in_cos113;
        8'b01110010 : cos2 = mux_in_cos114;
        8'b01110011 : cos2 = mux_in_cos115;
        8'b01110100 : cos2 = mux_in_cos116;
        8'b01110101 : cos2 = mux_in_cos117;
        8'b01110110 : cos2 = mux_in_cos118;
        8'b01110111 : cos2 = mux_in_cos119;
        8'b01111000 : cos2 = mux_in_cos120;
        8'b01111001 : cos2 = mux_in_cos121;
        8'b01111010 : cos2 = mux_in_cos122;
        8'b01111011 : cos2 = mux_in_cos123;
        8'b01111100 : cos2 = mux_in_cos124;
        8'b01111101 : cos2 = mux_in_cos125;
        8'b01111110 : cos2 = mux_in_cos126;
        8'b01111111 : cos2 = mux_in_cos127;
        8'b10000000 : cos2 = mux_in_cos128;
        default: cos2 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in3)
        8'b00000000 : cos3 = mux_in_cos0;
        8'b00000001 : cos3 = mux_in_cos1;
        8'b00000010 : cos3 = mux_in_cos2;
        8'b00000011 : cos3 = mux_in_cos3;
        8'b00000100 : cos3 = mux_in_cos4;
        8'b00000101 : cos3 = mux_in_cos5;
        8'b00000110 : cos3 = mux_in_cos6;
        8'b00000111 : cos3 = mux_in_cos7;
        8'b00001000 : cos3 = mux_in_cos8;
        8'b00001001 : cos3 = mux_in_cos9;
        8'b00001010 : cos3 = mux_in_cos10;
        8'b00001011 : cos3 = mux_in_cos11;
        8'b00001100 : cos3 = mux_in_cos12;
        8'b00001101 : cos3 = mux_in_cos13;
        8'b00001110 : cos3 = mux_in_cos14;
        8'b00001111 : cos3 = mux_in_cos15;
        8'b00010000 : cos3 = mux_in_cos16;
        8'b00010001 : cos3 = mux_in_cos17;
        8'b00010010 : cos3 = mux_in_cos18;
        8'b00010011 : cos3 = mux_in_cos19;
        8'b00010100 : cos3 = mux_in_cos20;
        8'b00010101 : cos3 = mux_in_cos21;
        8'b00010110 : cos3 = mux_in_cos22;
        8'b00010111 : cos3 = mux_in_cos23;
        8'b00011000 : cos3 = mux_in_cos24;
        8'b00011001 : cos3 = mux_in_cos25;
        8'b00011010 : cos3 = mux_in_cos26;
        8'b00011011 : cos3 = mux_in_cos27;
        8'b00011100 : cos3 = mux_in_cos28;
        8'b00011101 : cos3 = mux_in_cos29;
        8'b00011110 : cos3 = mux_in_cos30;
        8'b00011111 : cos3 = mux_in_cos31;
        8'b00100000 : cos3 = mux_in_cos32;
        8'b00100001 : cos3 = mux_in_cos33;
        8'b00100010 : cos3 = mux_in_cos34;
        8'b00100011 : cos3 = mux_in_cos35;
        8'b00100100 : cos3 = mux_in_cos36;
        8'b00100101 : cos3 = mux_in_cos37;
        8'b00100110 : cos3 = mux_in_cos38;
        8'b00100111 : cos3 = mux_in_cos39;
        8'b00101000 : cos3 = mux_in_cos40;
        8'b00101001 : cos3 = mux_in_cos41;
        8'b00101010 : cos3 = mux_in_cos42;
        8'b00101011 : cos3 = mux_in_cos43;
        8'b00101100 : cos3 = mux_in_cos44;
        8'b00101101 : cos3 = mux_in_cos45;
        8'b00101110 : cos3 = mux_in_cos46;
        8'b00101111 : cos3 = mux_in_cos47;
        8'b00110000 : cos3 = mux_in_cos48;
        8'b00110001 : cos3 = mux_in_cos49;
        8'b00110010 : cos3 = mux_in_cos50;
        8'b00110011 : cos3 = mux_in_cos51;
        8'b00110100 : cos3 = mux_in_cos52;
        8'b00110101 : cos3 = mux_in_cos53;
        8'b00110110 : cos3 = mux_in_cos54;
        8'b00110111 : cos3 = mux_in_cos55;
        8'b00111000 : cos3 = mux_in_cos56;
        8'b00111001 : cos3 = mux_in_cos57;
        8'b00111010 : cos3 = mux_in_cos58;
        8'b00111011 : cos3 = mux_in_cos59;
        8'b00111100 : cos3 = mux_in_cos60;
        8'b00111101 : cos3 = mux_in_cos61;
        8'b00111110 : cos3 = mux_in_cos62;
        8'b00111111 : cos3 = mux_in_cos63;
        8'b01000000 : cos3 = mux_in_cos64;
        8'b01000001 : cos3 = mux_in_cos65;
        8'b01000010 : cos3 = mux_in_cos66;
        8'b01000011 : cos3 = mux_in_cos67;
        8'b01000100 : cos3 = mux_in_cos68;
        8'b01000101 : cos3 = mux_in_cos69;
        8'b01000110 : cos3 = mux_in_cos70;
        8'b01000111 : cos3 = mux_in_cos71;
        8'b01001000 : cos3 = mux_in_cos72;
        8'b01001001 : cos3 = mux_in_cos73;
        8'b01001010 : cos3 = mux_in_cos74;
        8'b01001011 : cos3 = mux_in_cos75;
        8'b01001100 : cos3 = mux_in_cos76;
        8'b01001101 : cos3 = mux_in_cos77;
        8'b01001110 : cos3 = mux_in_cos78;
        8'b01001111 : cos3 = mux_in_cos79;
        8'b01010000 : cos3 = mux_in_cos80;
        8'b01010001 : cos3 = mux_in_cos81;
        8'b01010010 : cos3 = mux_in_cos82;
        8'b01010011 : cos3 = mux_in_cos83;
        8'b01010100 : cos3 = mux_in_cos84;
        8'b01010101 : cos3 = mux_in_cos85;
        8'b01010110 : cos3 = mux_in_cos86;
        8'b01010111 : cos3 = mux_in_cos87;
        8'b01011000 : cos3 = mux_in_cos88;
        8'b01011001 : cos3 = mux_in_cos89;
        8'b01011010 : cos3 = mux_in_cos90;
        8'b01011011 : cos3 = mux_in_cos91;
        8'b01011100 : cos3 = mux_in_cos92;
        8'b01011101 : cos3 = mux_in_cos93;
        8'b01011110 : cos3 = mux_in_cos94;
        8'b01011111 : cos3 = mux_in_cos95;
        8'b01100000 : cos3 = mux_in_cos96;
        8'b01100001 : cos3 = mux_in_cos97;
        8'b01100010 : cos3 = mux_in_cos98;
        8'b01100011 : cos3 = mux_in_cos99;
        8'b01100100 : cos3 = mux_in_cos100;
        8'b01100101 : cos3 = mux_in_cos101;
        8'b01100110 : cos3 = mux_in_cos102;
        8'b01100111 : cos3 = mux_in_cos103;
        8'b01101000 : cos3 = mux_in_cos104;
        8'b01101001 : cos3 = mux_in_cos105;
        8'b01101010 : cos3 = mux_in_cos106;
        8'b01101011 : cos3 = mux_in_cos107;
        8'b01101100 : cos3 = mux_in_cos108;
        8'b01101101 : cos3 = mux_in_cos109;
        8'b01101110 : cos3 = mux_in_cos110;
        8'b01101111 : cos3 = mux_in_cos111;
        8'b01110000 : cos3 = mux_in_cos112;
        8'b01110001 : cos3 = mux_in_cos113;
        8'b01110010 : cos3 = mux_in_cos114;
        8'b01110011 : cos3 = mux_in_cos115;
        8'b01110100 : cos3 = mux_in_cos116;
        8'b01110101 : cos3 = mux_in_cos117;
        8'b01110110 : cos3 = mux_in_cos118;
        8'b01110111 : cos3 = mux_in_cos119;
        8'b01111000 : cos3 = mux_in_cos120;
        8'b01111001 : cos3 = mux_in_cos121;
        8'b01111010 : cos3 = mux_in_cos122;
        8'b01111011 : cos3 = mux_in_cos123;
        8'b01111100 : cos3 = mux_in_cos124;
        8'b01111101 : cos3 = mux_in_cos125;
        8'b01111110 : cos3 = mux_in_cos126;
        8'b01111111 : cos3 = mux_in_cos127;
        8'b10000000 : cos3 = mux_in_cos128;
        default: cos3 = 15'bx;
        endcase
    end

endmodule