`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author: Pavan Kumar
// Create Date: 09-10-2024
// Module name: sin_cos_LUT_7QP_QORD3.v
//////////////////////////////////////////////////////////////////////////////////

module sin_cos_LUT_7QP_QORD3
(
    input      [ 6:0] x_in1,
    output reg [15:0] sin1, cos1
);

    wire [15:0] mux_in_cos0, mux_in_sin0, mux_in_cos1, mux_in_sin1, mux_in_cos2, mux_in_sin2, mux_in_cos3, mux_in_sin3, mux_in_cos4, mux_in_sin4, mux_in_cos5, mux_in_sin5, mux_in_cos6, mux_in_sin6, mux_in_cos7, mux_in_sin7, mux_in_cos8, mux_in_sin8, mux_in_cos9, mux_in_sin9, mux_in_cos10, mux_in_sin10, mux_in_cos11, mux_in_sin11, mux_in_cos12, mux_in_sin12, mux_in_cos13, mux_in_sin13, mux_in_cos14, mux_in_sin14, mux_in_cos15, mux_in_sin15, mux_in_cos16, mux_in_sin16, mux_in_cos17, mux_in_sin17, mux_in_cos18, mux_in_sin18, mux_in_cos19, mux_in_sin19, mux_in_cos20, mux_in_sin20, mux_in_cos21, mux_in_sin21, mux_in_cos22, mux_in_sin22, mux_in_cos23, mux_in_sin23, mux_in_cos24, mux_in_sin24, mux_in_cos25, mux_in_sin25, mux_in_cos26, mux_in_sin26, mux_in_cos27, mux_in_sin27, mux_in_cos28, mux_in_sin28, mux_in_cos29, mux_in_sin29, mux_in_cos30, mux_in_sin30, mux_in_cos31, mux_in_sin31, mux_in_cos32, mux_in_sin32, mux_in_cos33, mux_in_sin33, mux_in_cos34, mux_in_sin34, mux_in_cos35, mux_in_sin35, mux_in_cos36, mux_in_sin36, mux_in_cos37, mux_in_sin37, mux_in_cos38, mux_in_sin38, mux_in_cos39, mux_in_sin39, mux_in_cos40, mux_in_sin40, mux_in_cos41, mux_in_sin41, mux_in_cos42, mux_in_sin42, mux_in_cos43, mux_in_sin43, mux_in_cos44, mux_in_sin44, mux_in_cos45, mux_in_sin45, mux_in_cos46, mux_in_sin46, mux_in_cos47, mux_in_sin47, mux_in_cos48, mux_in_sin48, mux_in_cos49, mux_in_sin49, mux_in_cos50, mux_in_sin50, mux_in_cos51, mux_in_sin51, mux_in_cos52, mux_in_sin52, mux_in_cos53, mux_in_sin53, mux_in_cos54, mux_in_sin54, mux_in_cos55, mux_in_sin55, mux_in_cos56, mux_in_sin56, mux_in_cos57, mux_in_sin57, mux_in_cos58, mux_in_sin58, mux_in_cos59, mux_in_sin59, mux_in_cos60, mux_in_sin60, mux_in_cos61, mux_in_sin61, mux_in_cos62, mux_in_sin62, mux_in_cos63, mux_in_sin63, mux_in_cos64, mux_in_sin64;

    assign mux_in_cos0 = 16'b1000000000000000;
    assign mux_in_sin0 = 16'b0000000000000000;
    assign mux_in_cos1 = 16'b0111111111110110;
    assign mux_in_sin1 = 16'b0000001100100100;
    assign mux_in_cos2 = 16'b0111111111011001;
    assign mux_in_sin2 = 16'b0000011001001000;
    assign mux_in_cos3 = 16'b0111111110100111;
    assign mux_in_sin3 = 16'b0000100101101011;
    assign mux_in_cos4 = 16'b0111111101100010;
    assign mux_in_sin4 = 16'b0000110010001100;
    assign mux_in_cos5 = 16'b0111111100001010;
    assign mux_in_sin5 = 16'b0000111110101011;
    assign mux_in_cos6 = 16'b0111111010011101;
    assign mux_in_sin6 = 16'b0001001011001000;
    assign mux_in_cos7 = 16'b0111111000011110;
    assign mux_in_sin7 = 16'b0001010111100010;
    assign mux_in_cos8 = 16'b0111110110001010;
    assign mux_in_sin8 = 16'b0001100011111001;
    assign mux_in_cos9 = 16'b0111110011100100;
    assign mux_in_sin9 = 16'b0001110000001100;
    assign mux_in_cos10 = 16'b0111110000101010;
    assign mux_in_sin10 = 16'b0001111100011010;
    assign mux_in_cos11 = 16'b0111101101011101;
    assign mux_in_sin11 = 16'b0010001000100100;
    assign mux_in_cos12 = 16'b0111101001111101;
    assign mux_in_sin12 = 16'b0010010100101000;
    assign mux_in_cos13 = 16'b0111100110001010;
    assign mux_in_sin13 = 16'b0010100000100111;
    assign mux_in_cos14 = 16'b0111100010000101;
    assign mux_in_sin14 = 16'b0010101100011111;
    assign mux_in_cos15 = 16'b0111011101101100;
    assign mux_in_sin15 = 16'b0010111000010001;
    assign mux_in_cos16 = 16'b0111011001000010;
    assign mux_in_sin16 = 16'b0011000011111100;
    assign mux_in_cos17 = 16'b0111010100000101;
    assign mux_in_sin17 = 16'b0011001111011111;
    assign mux_in_cos18 = 16'b0111001110110110;
    assign mux_in_sin18 = 16'b0011011010111010;
    assign mux_in_cos19 = 16'b0111001001010101;
    assign mux_in_sin19 = 16'b0011100110001101;
    assign mux_in_cos20 = 16'b0111000011100011;
    assign mux_in_sin20 = 16'b0011110001010111;
    assign mux_in_cos21 = 16'b0110111101011111;
    assign mux_in_sin21 = 16'b0011111100010111;
    assign mux_in_cos22 = 16'b0110110111001010;
    assign mux_in_sin22 = 16'b0100000111001110;
    assign mux_in_cos23 = 16'b0110110000100100;
    assign mux_in_sin23 = 16'b0100010001111011;
    assign mux_in_cos24 = 16'b0110101001101110;
    assign mux_in_sin24 = 16'b0100011100011101;
    assign mux_in_cos25 = 16'b0110100010100111;
    assign mux_in_sin25 = 16'b0100100110110100;
    assign mux_in_cos26 = 16'b0110011011010000;
    assign mux_in_sin26 = 16'b0100110001000000;
    assign mux_in_cos27 = 16'b0110010011101001;
    assign mux_in_sin27 = 16'b0100111011000000;
    assign mux_in_cos28 = 16'b0110001011110010;
    assign mux_in_sin28 = 16'b0101000100110100;
    assign mux_in_cos29 = 16'b0110000011101100;
    assign mux_in_sin29 = 16'b0101001110011011;
    assign mux_in_cos30 = 16'b0101111011010111;
    assign mux_in_sin30 = 16'b0101010111110110;
    assign mux_in_cos31 = 16'b0101110010110100;
    assign mux_in_sin31 = 16'b0101100001000011;
    assign mux_in_cos32 = 16'b0101101010000010;
    assign mux_in_sin32 = 16'b0101101010000010;
    assign mux_in_cos33 = 16'b0101100001000011;
    assign mux_in_sin33 = 16'b0101110010110100;
    assign mux_in_cos34 = 16'b0101010111110110;
    assign mux_in_sin34 = 16'b0101111011010111;
    assign mux_in_cos35 = 16'b0101001110011011;
    assign mux_in_sin35 = 16'b0110000011101100;
    assign mux_in_cos36 = 16'b0101000100110100;
    assign mux_in_sin36 = 16'b0110001011110010;
    assign mux_in_cos37 = 16'b0100111011000000;
    assign mux_in_sin37 = 16'b0110010011101001;
    assign mux_in_cos38 = 16'b0100110001000000;
    assign mux_in_sin38 = 16'b0110011011010000;
    assign mux_in_cos39 = 16'b0100100110110100;
    assign mux_in_sin39 = 16'b0110100010100111;
    assign mux_in_cos40 = 16'b0100011100011101;
    assign mux_in_sin40 = 16'b0110101001101110;
    assign mux_in_cos41 = 16'b0100010001111011;
    assign mux_in_sin41 = 16'b0110110000100100;
    assign mux_in_cos42 = 16'b0100000111001110;
    assign mux_in_sin42 = 16'b0110110111001010;
    assign mux_in_cos43 = 16'b0011111100010111;
    assign mux_in_sin43 = 16'b0110111101011111;
    assign mux_in_cos44 = 16'b0011110001010111;
    assign mux_in_sin44 = 16'b0111000011100011;
    assign mux_in_cos45 = 16'b0011100110001101;
    assign mux_in_sin45 = 16'b0111001001010101;
    assign mux_in_cos46 = 16'b0011011010111010;
    assign mux_in_sin46 = 16'b0111001110110110;
    assign mux_in_cos47 = 16'b0011001111011111;
    assign mux_in_sin47 = 16'b0111010100000101;
    assign mux_in_cos48 = 16'b0011000011111100;
    assign mux_in_sin48 = 16'b0111011001000010;
    assign mux_in_cos49 = 16'b0010111000010001;
    assign mux_in_sin49 = 16'b0111011101101100;
    assign mux_in_cos50 = 16'b0010101100011111;
    assign mux_in_sin50 = 16'b0111100010000101;
    assign mux_in_cos51 = 16'b0010100000100111;
    assign mux_in_sin51 = 16'b0111100110001010;
    assign mux_in_cos52 = 16'b0010010100101000;
    assign mux_in_sin52 = 16'b0111101001111101;
    assign mux_in_cos53 = 16'b0010001000100100;
    assign mux_in_sin53 = 16'b0111101101011101;
    assign mux_in_cos54 = 16'b0001111100011010;
    assign mux_in_sin54 = 16'b0111110000101010;
    assign mux_in_cos55 = 16'b0001110000001100;
    assign mux_in_sin55 = 16'b0111110011100100;
    assign mux_in_cos56 = 16'b0001100011111001;
    assign mux_in_sin56 = 16'b0111110110001010;
    assign mux_in_cos57 = 16'b0001010111100010;
    assign mux_in_sin57 = 16'b0111111000011110;
    assign mux_in_cos58 = 16'b0001001011001000;
    assign mux_in_sin58 = 16'b0111111010011101;
    assign mux_in_cos59 = 16'b0000111110101011;
    assign mux_in_sin59 = 16'b0111111100001010;
    assign mux_in_cos60 = 16'b0000110010001100;
    assign mux_in_sin60 = 16'b0111111101100010;
    assign mux_in_cos61 = 16'b0000100101101011;
    assign mux_in_sin61 = 16'b0111111110100111;
    assign mux_in_cos62 = 16'b0000011001001000;
    assign mux_in_sin62 = 16'b0111111111011001;
    assign mux_in_cos63 = 16'b0000001100100100;
    assign mux_in_sin63 = 16'b0111111111110110;
    assign mux_in_cos64 = 16'b0000000000000000;
    assign mux_in_sin64 = 16'b1000000000000000;

    // Sine LUTs

    always @ (*)
    begin
        case(x_in1)
        7'b0000000 : sin1 = mux_in_sin0;
        7'b0000001 : sin1 = mux_in_sin1;
        7'b0000010 : sin1 = mux_in_sin2;
        7'b0000011 : sin1 = mux_in_sin3;
        7'b0000100 : sin1 = mux_in_sin4;
        7'b0000101 : sin1 = mux_in_sin5;
        7'b0000110 : sin1 = mux_in_sin6;
        7'b0000111 : sin1 = mux_in_sin7;
        7'b0001000 : sin1 = mux_in_sin8;
        7'b0001001 : sin1 = mux_in_sin9;
        7'b0001010 : sin1 = mux_in_sin10;
        7'b0001011 : sin1 = mux_in_sin11;
        7'b0001100 : sin1 = mux_in_sin12;
        7'b0001101 : sin1 = mux_in_sin13;
        7'b0001110 : sin1 = mux_in_sin14;
        7'b0001111 : sin1 = mux_in_sin15;
        7'b0010000 : sin1 = mux_in_sin16;
        7'b0010001 : sin1 = mux_in_sin17;
        7'b0010010 : sin1 = mux_in_sin18;
        7'b0010011 : sin1 = mux_in_sin19;
        7'b0010100 : sin1 = mux_in_sin20;
        7'b0010101 : sin1 = mux_in_sin21;
        7'b0010110 : sin1 = mux_in_sin22;
        7'b0010111 : sin1 = mux_in_sin23;
        7'b0011000 : sin1 = mux_in_sin24;
        7'b0011001 : sin1 = mux_in_sin25;
        7'b0011010 : sin1 = mux_in_sin26;
        7'b0011011 : sin1 = mux_in_sin27;
        7'b0011100 : sin1 = mux_in_sin28;
        7'b0011101 : sin1 = mux_in_sin29;
        7'b0011110 : sin1 = mux_in_sin30;
        7'b0011111 : sin1 = mux_in_sin31;
        7'b0100000 : sin1 = mux_in_sin32;
        7'b0100001 : sin1 = mux_in_sin33;
        7'b0100010 : sin1 = mux_in_sin34;
        7'b0100011 : sin1 = mux_in_sin35;
        7'b0100100 : sin1 = mux_in_sin36;
        7'b0100101 : sin1 = mux_in_sin37;
        7'b0100110 : sin1 = mux_in_sin38;
        7'b0100111 : sin1 = mux_in_sin39;
        7'b0101000 : sin1 = mux_in_sin40;
        7'b0101001 : sin1 = mux_in_sin41;
        7'b0101010 : sin1 = mux_in_sin42;
        7'b0101011 : sin1 = mux_in_sin43;
        7'b0101100 : sin1 = mux_in_sin44;
        7'b0101101 : sin1 = mux_in_sin45;
        7'b0101110 : sin1 = mux_in_sin46;
        7'b0101111 : sin1 = mux_in_sin47;
        7'b0110000 : sin1 = mux_in_sin48;
        7'b0110001 : sin1 = mux_in_sin49;
        7'b0110010 : sin1 = mux_in_sin50;
        7'b0110011 : sin1 = mux_in_sin51;
        7'b0110100 : sin1 = mux_in_sin52;
        7'b0110101 : sin1 = mux_in_sin53;
        7'b0110110 : sin1 = mux_in_sin54;
        7'b0110111 : sin1 = mux_in_sin55;
        7'b0111000 : sin1 = mux_in_sin56;
        7'b0111001 : sin1 = mux_in_sin57;
        7'b0111010 : sin1 = mux_in_sin58;
        7'b0111011 : sin1 = mux_in_sin59;
        7'b0111100 : sin1 = mux_in_sin60;
        7'b0111101 : sin1 = mux_in_sin61;
        7'b0111110 : sin1 = mux_in_sin62;
        7'b0111111 : sin1 = mux_in_sin63;
        7'b1000000 : sin1 = mux_in_sin64;
        default: sin1 = 15'bx;
        endcase
    end

    //Cos LUTs
    always @ (*)
    begin
        case(x_in1)
        7'b0000000 : cos1 = mux_in_cos0;
        7'b0000001 : cos1 = mux_in_cos1;
        7'b0000010 : cos1 = mux_in_cos2;
        7'b0000011 : cos1 = mux_in_cos3;
        7'b0000100 : cos1 = mux_in_cos4;
        7'b0000101 : cos1 = mux_in_cos5;
        7'b0000110 : cos1 = mux_in_cos6;
        7'b0000111 : cos1 = mux_in_cos7;
        7'b0001000 : cos1 = mux_in_cos8;
        7'b0001001 : cos1 = mux_in_cos9;
        7'b0001010 : cos1 = mux_in_cos10;
        7'b0001011 : cos1 = mux_in_cos11;
        7'b0001100 : cos1 = mux_in_cos12;
        7'b0001101 : cos1 = mux_in_cos13;
        7'b0001110 : cos1 = mux_in_cos14;
        7'b0001111 : cos1 = mux_in_cos15;
        7'b0010000 : cos1 = mux_in_cos16;
        7'b0010001 : cos1 = mux_in_cos17;
        7'b0010010 : cos1 = mux_in_cos18;
        7'b0010011 : cos1 = mux_in_cos19;
        7'b0010100 : cos1 = mux_in_cos20;
        7'b0010101 : cos1 = mux_in_cos21;
        7'b0010110 : cos1 = mux_in_cos22;
        7'b0010111 : cos1 = mux_in_cos23;
        7'b0011000 : cos1 = mux_in_cos24;
        7'b0011001 : cos1 = mux_in_cos25;
        7'b0011010 : cos1 = mux_in_cos26;
        7'b0011011 : cos1 = mux_in_cos27;
        7'b0011100 : cos1 = mux_in_cos28;
        7'b0011101 : cos1 = mux_in_cos29;
        7'b0011110 : cos1 = mux_in_cos30;
        7'b0011111 : cos1 = mux_in_cos31;
        7'b0100000 : cos1 = mux_in_cos32;
        7'b0100001 : cos1 = mux_in_cos33;
        7'b0100010 : cos1 = mux_in_cos34;
        7'b0100011 : cos1 = mux_in_cos35;
        7'b0100100 : cos1 = mux_in_cos36;
        7'b0100101 : cos1 = mux_in_cos37;
        7'b0100110 : cos1 = mux_in_cos38;
        7'b0100111 : cos1 = mux_in_cos39;
        7'b0101000 : cos1 = mux_in_cos40;
        7'b0101001 : cos1 = mux_in_cos41;
        7'b0101010 : cos1 = mux_in_cos42;
        7'b0101011 : cos1 = mux_in_cos43;
        7'b0101100 : cos1 = mux_in_cos44;
        7'b0101101 : cos1 = mux_in_cos45;
        7'b0101110 : cos1 = mux_in_cos46;
        7'b0101111 : cos1 = mux_in_cos47;
        7'b0110000 : cos1 = mux_in_cos48;
        7'b0110001 : cos1 = mux_in_cos49;
        7'b0110010 : cos1 = mux_in_cos50;
        7'b0110011 : cos1 = mux_in_cos51;
        7'b0110100 : cos1 = mux_in_cos52;
        7'b0110101 : cos1 = mux_in_cos53;
        7'b0110110 : cos1 = mux_in_cos54;
        7'b0110111 : cos1 = mux_in_cos55;
        7'b0111000 : cos1 = mux_in_cos56;
        7'b0111001 : cos1 = mux_in_cos57;
        7'b0111010 : cos1 = mux_in_cos58;
        7'b0111011 : cos1 = mux_in_cos59;
        7'b0111100 : cos1 = mux_in_cos60;
        7'b0111101 : cos1 = mux_in_cos61;
        7'b0111110 : cos1 = mux_in_cos62;
        7'b0111111 : cos1 = mux_in_cos63;
        7'b1000000 : cos1 = mux_in_cos64;
        default: cos1 = 15'bx;
        endcase
    end


endmodule