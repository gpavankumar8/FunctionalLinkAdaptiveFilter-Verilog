`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author: Pavan Kumar
// Create Date: 29-07-2024
// Module name: log_sin_cos_LUT_9QP.v
//////////////////////////////////////////////////////////////////////////////////

module log_sin_cos_LUT_9QP
(
    input      [ 8:0] x_in1, x_in2, x_in3,
    output reg [15:0] logsin1, logsin2, logsin3, logcos1, logcos2, logcos3
);

    wire [15:0] mux_in_cos0, mux_in_sin0, mux_in_cos1, mux_in_sin1, mux_in_cos2, mux_in_sin2, mux_in_cos3, mux_in_sin3, mux_in_cos4, mux_in_sin4, mux_in_cos5, mux_in_sin5, mux_in_cos6, mux_in_sin6, mux_in_cos7, mux_in_sin7, mux_in_cos8, mux_in_sin8, mux_in_cos9, mux_in_sin9, mux_in_cos10, mux_in_sin10, mux_in_cos11, mux_in_sin11, mux_in_cos12, mux_in_sin12, mux_in_cos13, mux_in_sin13, mux_in_cos14, mux_in_sin14, mux_in_cos15, mux_in_sin15, mux_in_cos16, mux_in_sin16, mux_in_cos17, mux_in_sin17, mux_in_cos18, mux_in_sin18, mux_in_cos19, mux_in_sin19, mux_in_cos20, mux_in_sin20, mux_in_cos21, mux_in_sin21, mux_in_cos22, mux_in_sin22, mux_in_cos23, mux_in_sin23, mux_in_cos24, mux_in_sin24, mux_in_cos25, mux_in_sin25, mux_in_cos26, mux_in_sin26, mux_in_cos27, mux_in_sin27, mux_in_cos28, mux_in_sin28, mux_in_cos29, mux_in_sin29, mux_in_cos30, mux_in_sin30, mux_in_cos31, mux_in_sin31, mux_in_cos32, mux_in_sin32, mux_in_cos33, mux_in_sin33, mux_in_cos34, mux_in_sin34, mux_in_cos35, mux_in_sin35, mux_in_cos36, mux_in_sin36, mux_in_cos37, mux_in_sin37, mux_in_cos38, mux_in_sin38, mux_in_cos39, mux_in_sin39, mux_in_cos40, mux_in_sin40, mux_in_cos41, mux_in_sin41, mux_in_cos42, mux_in_sin42, mux_in_cos43, mux_in_sin43, mux_in_cos44, mux_in_sin44, mux_in_cos45, mux_in_sin45, mux_in_cos46, mux_in_sin46, mux_in_cos47, mux_in_sin47, mux_in_cos48, mux_in_sin48, mux_in_cos49, mux_in_sin49, mux_in_cos50, mux_in_sin50, mux_in_cos51, mux_in_sin51, mux_in_cos52, mux_in_sin52, mux_in_cos53, mux_in_sin53, mux_in_cos54, mux_in_sin54, mux_in_cos55, mux_in_sin55, mux_in_cos56, mux_in_sin56, mux_in_cos57, mux_in_sin57, mux_in_cos58, mux_in_sin58, mux_in_cos59, mux_in_sin59, mux_in_cos60, mux_in_sin60, mux_in_cos61, mux_in_sin61, mux_in_cos62, mux_in_sin62, mux_in_cos63, mux_in_sin63, mux_in_cos64, mux_in_sin64, mux_in_cos65, mux_in_sin65, mux_in_cos66, mux_in_sin66, mux_in_cos67, mux_in_sin67, mux_in_cos68, mux_in_sin68, mux_in_cos69, mux_in_sin69, mux_in_cos70, mux_in_sin70, mux_in_cos71, mux_in_sin71, mux_in_cos72, mux_in_sin72, mux_in_cos73, mux_in_sin73, mux_in_cos74, mux_in_sin74, mux_in_cos75, mux_in_sin75, mux_in_cos76, mux_in_sin76, mux_in_cos77, mux_in_sin77, mux_in_cos78, mux_in_sin78, mux_in_cos79, mux_in_sin79, mux_in_cos80, mux_in_sin80, mux_in_cos81, mux_in_sin81, mux_in_cos82, mux_in_sin82, mux_in_cos83, mux_in_sin83, mux_in_cos84, mux_in_sin84, mux_in_cos85, mux_in_sin85, mux_in_cos86, mux_in_sin86, mux_in_cos87, mux_in_sin87, mux_in_cos88, mux_in_sin88, mux_in_cos89, mux_in_sin89, mux_in_cos90, mux_in_sin90, mux_in_cos91, mux_in_sin91, mux_in_cos92, mux_in_sin92, mux_in_cos93, mux_in_sin93, mux_in_cos94, mux_in_sin94, mux_in_cos95, mux_in_sin95, mux_in_cos96, mux_in_sin96, mux_in_cos97, mux_in_sin97, mux_in_cos98, mux_in_sin98, mux_in_cos99, mux_in_sin99, mux_in_cos100, mux_in_sin100, mux_in_cos101, mux_in_sin101, mux_in_cos102, mux_in_sin102, mux_in_cos103, mux_in_sin103, mux_in_cos104, mux_in_sin104, mux_in_cos105, mux_in_sin105, mux_in_cos106, mux_in_sin106, mux_in_cos107, mux_in_sin107, mux_in_cos108, mux_in_sin108, mux_in_cos109, mux_in_sin109, mux_in_cos110, mux_in_sin110, mux_in_cos111, mux_in_sin111, mux_in_cos112, mux_in_sin112, mux_in_cos113, mux_in_sin113, mux_in_cos114, mux_in_sin114, mux_in_cos115, mux_in_sin115, mux_in_cos116, mux_in_sin116, mux_in_cos117, mux_in_sin117, mux_in_cos118, mux_in_sin118, mux_in_cos119, mux_in_sin119, mux_in_cos120, mux_in_sin120, mux_in_cos121, mux_in_sin121, mux_in_cos122, mux_in_sin122, mux_in_cos123, mux_in_sin123, mux_in_cos124, mux_in_sin124, mux_in_cos125, mux_in_sin125, mux_in_cos126, mux_in_sin126, mux_in_cos127, mux_in_sin127, mux_in_cos128, mux_in_sin128, mux_in_cos129, mux_in_sin129, mux_in_cos130, mux_in_sin130, mux_in_cos131, mux_in_sin131, mux_in_cos132, mux_in_sin132, mux_in_cos133, mux_in_sin133, mux_in_cos134, mux_in_sin134, mux_in_cos135, mux_in_sin135, mux_in_cos136, mux_in_sin136, mux_in_cos137, mux_in_sin137, mux_in_cos138, mux_in_sin138, mux_in_cos139, mux_in_sin139, mux_in_cos140, mux_in_sin140, mux_in_cos141, mux_in_sin141, mux_in_cos142, mux_in_sin142, mux_in_cos143, mux_in_sin143, mux_in_cos144, mux_in_sin144, mux_in_cos145, mux_in_sin145, mux_in_cos146, mux_in_sin146, mux_in_cos147, mux_in_sin147, mux_in_cos148, mux_in_sin148, mux_in_cos149, mux_in_sin149, mux_in_cos150, mux_in_sin150, mux_in_cos151, mux_in_sin151, mux_in_cos152, mux_in_sin152, mux_in_cos153, mux_in_sin153, mux_in_cos154, mux_in_sin154, mux_in_cos155, mux_in_sin155, mux_in_cos156, mux_in_sin156, mux_in_cos157, mux_in_sin157, mux_in_cos158, mux_in_sin158, mux_in_cos159, mux_in_sin159, mux_in_cos160, mux_in_sin160, mux_in_cos161, mux_in_sin161, mux_in_cos162, mux_in_sin162, mux_in_cos163, mux_in_sin163, mux_in_cos164, mux_in_sin164, mux_in_cos165, mux_in_sin165, mux_in_cos166, mux_in_sin166, mux_in_cos167, mux_in_sin167, mux_in_cos168, mux_in_sin168, mux_in_cos169, mux_in_sin169, mux_in_cos170, mux_in_sin170, mux_in_cos171, mux_in_sin171, mux_in_cos172, mux_in_sin172, mux_in_cos173, mux_in_sin173, mux_in_cos174, mux_in_sin174, mux_in_cos175, mux_in_sin175, mux_in_cos176, mux_in_sin176, mux_in_cos177, mux_in_sin177, mux_in_cos178, mux_in_sin178, mux_in_cos179, mux_in_sin179, mux_in_cos180, mux_in_sin180, mux_in_cos181, mux_in_sin181, mux_in_cos182, mux_in_sin182, mux_in_cos183, mux_in_sin183, mux_in_cos184, mux_in_sin184, mux_in_cos185, mux_in_sin185, mux_in_cos186, mux_in_sin186, mux_in_cos187, mux_in_sin187, mux_in_cos188, mux_in_sin188, mux_in_cos189, mux_in_sin189, mux_in_cos190, mux_in_sin190, mux_in_cos191, mux_in_sin191, mux_in_cos192, mux_in_sin192, mux_in_cos193, mux_in_sin193, mux_in_cos194, mux_in_sin194, mux_in_cos195, mux_in_sin195, mux_in_cos196, mux_in_sin196, mux_in_cos197, mux_in_sin197, mux_in_cos198, mux_in_sin198, mux_in_cos199, mux_in_sin199, mux_in_cos200, mux_in_sin200, mux_in_cos201, mux_in_sin201, mux_in_cos202, mux_in_sin202, mux_in_cos203, mux_in_sin203, mux_in_cos204, mux_in_sin204, mux_in_cos205, mux_in_sin205, mux_in_cos206, mux_in_sin206, mux_in_cos207, mux_in_sin207, mux_in_cos208, mux_in_sin208, mux_in_cos209, mux_in_sin209, mux_in_cos210, mux_in_sin210, mux_in_cos211, mux_in_sin211, mux_in_cos212, mux_in_sin212, mux_in_cos213, mux_in_sin213, mux_in_cos214, mux_in_sin214, mux_in_cos215, mux_in_sin215, mux_in_cos216, mux_in_sin216, mux_in_cos217, mux_in_sin217, mux_in_cos218, mux_in_sin218, mux_in_cos219, mux_in_sin219, mux_in_cos220, mux_in_sin220, mux_in_cos221, mux_in_sin221, mux_in_cos222, mux_in_sin222, mux_in_cos223, mux_in_sin223, mux_in_cos224, mux_in_sin224, mux_in_cos225, mux_in_sin225, mux_in_cos226, mux_in_sin226, mux_in_cos227, mux_in_sin227, mux_in_cos228, mux_in_sin228, mux_in_cos229, mux_in_sin229, mux_in_cos230, mux_in_sin230, mux_in_cos231, mux_in_sin231, mux_in_cos232, mux_in_sin232, mux_in_cos233, mux_in_sin233, mux_in_cos234, mux_in_sin234, mux_in_cos235, mux_in_sin235, mux_in_cos236, mux_in_sin236, mux_in_cos237, mux_in_sin237, mux_in_cos238, mux_in_sin238, mux_in_cos239, mux_in_sin239, mux_in_cos240, mux_in_sin240, mux_in_cos241, mux_in_sin241, mux_in_cos242, mux_in_sin242, mux_in_cos243, mux_in_sin243, mux_in_cos244, mux_in_sin244, mux_in_cos245, mux_in_sin245, mux_in_cos246, mux_in_sin246, mux_in_cos247, mux_in_sin247, mux_in_cos248, mux_in_sin248, mux_in_cos249, mux_in_sin249, mux_in_cos250, mux_in_sin250, mux_in_cos251, mux_in_sin251, mux_in_cos252, mux_in_sin252, mux_in_cos253, mux_in_sin253, mux_in_cos254, mux_in_sin254, mux_in_cos255, mux_in_sin255, mux_in_cos256, mux_in_sin256;

    assign mux_in_cos0 = 16'b0000000000000000;
    assign mux_in_sin0 = 16'b0000000000000000;
    assign mux_in_cos1 = 16'b0000000000000000;
    assign mux_in_sin1 = 16'b1000101001101100;
    assign mux_in_cos2 = 16'b0000000000000000;
    assign mux_in_sin2 = 16'b1001101001101100;
    assign mux_in_cos3 = 16'b1111111111111111;
    assign mux_in_sin3 = 16'b1010001111001000;
    assign mux_in_cos4 = 16'b1111111111111110;
    assign mux_in_sin4 = 16'b1010101001101100;
    assign mux_in_cos5 = 16'b1111111111111101;
    assign mux_in_sin5 = 16'b1010111110010010;
    assign mux_in_cos6 = 16'b1111111111111100;
    assign mux_in_sin6 = 16'b1011001111000111;
    assign mux_in_cos7 = 16'b1111111111111011;
    assign mux_in_sin7 = 16'b1011011101010110;
    assign mux_in_cos8 = 16'b1111111111111001;
    assign mux_in_sin8 = 16'b1011101001101010;
    assign mux_in_cos9 = 16'b1111111111110111;
    assign mux_in_sin9 = 16'b1011110100100010;
    assign mux_in_cos10 = 16'b1111111111110101;
    assign mux_in_sin10 = 16'b1011111110001111;
    assign mux_in_cos11 = 16'b1111111111110011;
    assign mux_in_sin11 = 16'b1100000111000010;
    assign mux_in_cos12 = 16'b1111111111110000;
    assign mux_in_sin12 = 16'b1100001111000011;
    assign mux_in_cos13 = 16'b1111111111101101;
    assign mux_in_sin13 = 16'b1100010110011011;
    assign mux_in_cos14 = 16'b1111111111101010;
    assign mux_in_sin14 = 16'b1100011101010000;
    assign mux_in_cos15 = 16'b1111111111100111;
    assign mux_in_sin15 = 16'b1100100011100111;
    assign mux_in_cos16 = 16'b1111111111100011;
    assign mux_in_sin16 = 16'b1100101001100011;
    assign mux_in_cos17 = 16'b1111111111100000;
    assign mux_in_sin17 = 16'b1100101111001000;
    assign mux_in_cos18 = 16'b1111111111011100;
    assign mux_in_sin18 = 16'b1100110100011001;
    assign mux_in_cos19 = 16'b1111111111011000;
    assign mux_in_sin19 = 16'b1100111001010111;
    assign mux_in_cos20 = 16'b1111111111010011;
    assign mux_in_sin20 = 16'b1100111110000100;
    assign mux_in_cos21 = 16'b1111111111001111;
    assign mux_in_sin21 = 16'b1101000010100011;
    assign mux_in_cos22 = 16'b1111111111001010;
    assign mux_in_sin22 = 16'b1101000110110100;
    assign mux_in_cos23 = 16'b1111111111000101;
    assign mux_in_sin23 = 16'b1101001010111001;
    assign mux_in_cos24 = 16'b1111111111000000;
    assign mux_in_sin24 = 16'b1101001110110011;
    assign mux_in_cos25 = 16'b1111111110111010;
    assign mux_in_sin25 = 16'b1101010010100011;
    assign mux_in_cos26 = 16'b1111111110110100;
    assign mux_in_sin26 = 16'b1101010110001000;
    assign mux_in_cos27 = 16'b1111111110101111;
    assign mux_in_sin27 = 16'b1101011001100101;
    assign mux_in_cos28 = 16'b1111111110101000;
    assign mux_in_sin28 = 16'b1101011100111010;
    assign mux_in_cos29 = 16'b1111111110100010;
    assign mux_in_sin29 = 16'b1101100000001000;
    assign mux_in_cos30 = 16'b1111111110011011;
    assign mux_in_sin30 = 16'b1101100011001110;
    assign mux_in_cos31 = 16'b1111111110010100;
    assign mux_in_sin31 = 16'b1101100110001101;
    assign mux_in_cos32 = 16'b1111111110001101;
    assign mux_in_sin32 = 16'b1101101001000111;
    assign mux_in_cos33 = 16'b1111111110000110;
    assign mux_in_sin33 = 16'b1101101011111010;
    assign mux_in_cos34 = 16'b1111111101111110;
    assign mux_in_sin34 = 16'b1101101110101000;
    assign mux_in_cos35 = 16'b1111111101110111;
    assign mux_in_sin35 = 16'b1101110001010001;
    assign mux_in_cos36 = 16'b1111111101101111;
    assign mux_in_sin36 = 16'b1101110011110100;
    assign mux_in_cos37 = 16'b1111111101100110;
    assign mux_in_sin37 = 16'b1101110110010100;
    assign mux_in_cos38 = 16'b1111111101011110;
    assign mux_in_sin38 = 16'b1101111000101110;
    assign mux_in_cos39 = 16'b1111111101010101;
    assign mux_in_sin39 = 16'b1101111011000101;
    assign mux_in_cos40 = 16'b1111111101001100;
    assign mux_in_sin40 = 16'b1101111101011000;
    assign mux_in_cos41 = 16'b1111111101000011;
    assign mux_in_sin41 = 16'b1101111111100111;
    assign mux_in_cos42 = 16'b1111111100111010;
    assign mux_in_sin42 = 16'b1110000001110010;
    assign mux_in_cos43 = 16'b1111111100110000;
    assign mux_in_sin43 = 16'b1110000011111010;
    assign mux_in_cos44 = 16'b1111111100100110;
    assign mux_in_sin44 = 16'b1110000101111110;
    assign mux_in_cos45 = 16'b1111111100011100;
    assign mux_in_sin45 = 16'b1110001000000000;
    assign mux_in_cos46 = 16'b1111111100010001;
    assign mux_in_sin46 = 16'b1110001001111110;
    assign mux_in_cos47 = 16'b1111111100000111;
    assign mux_in_sin47 = 16'b1110001011111010;
    assign mux_in_cos48 = 16'b1111111011111100;
    assign mux_in_sin48 = 16'b1110001101110011;
    assign mux_in_cos49 = 16'b1111111011110001;
    assign mux_in_sin49 = 16'b1110001111101001;
    assign mux_in_cos50 = 16'b1111111011100101;
    assign mux_in_sin50 = 16'b1110010001011101;
    assign mux_in_cos51 = 16'b1111111011011010;
    assign mux_in_sin51 = 16'b1110010011001110;
    assign mux_in_cos52 = 16'b1111111011001110;
    assign mux_in_sin52 = 16'b1110010100111101;
    assign mux_in_cos53 = 16'b1111111011000010;
    assign mux_in_sin53 = 16'b1110010110101010;
    assign mux_in_cos54 = 16'b1111111010110110;
    assign mux_in_sin54 = 16'b1110011000010100;
    assign mux_in_cos55 = 16'b1111111010101001;
    assign mux_in_sin55 = 16'b1110011001111100;
    assign mux_in_cos56 = 16'b1111111010011100;
    assign mux_in_sin56 = 16'b1110011011100011;
    assign mux_in_cos57 = 16'b1111111010001111;
    assign mux_in_sin57 = 16'b1110011101000111;
    assign mux_in_cos58 = 16'b1111111010000010;
    assign mux_in_sin58 = 16'b1110011110101010;
    assign mux_in_cos59 = 16'b1111111001110100;
    assign mux_in_sin59 = 16'b1110100000001010;
    assign mux_in_cos60 = 16'b1111111001100110;
    assign mux_in_sin60 = 16'b1110100001101001;
    assign mux_in_cos61 = 16'b1111111001011000;
    assign mux_in_sin61 = 16'b1110100011000110;
    assign mux_in_cos62 = 16'b1111111001001010;
    assign mux_in_sin62 = 16'b1110100100100010;
    assign mux_in_cos63 = 16'b1111111000111011;
    assign mux_in_sin63 = 16'b1110100101111100;
    assign mux_in_cos64 = 16'b1111111000101100;
    assign mux_in_sin64 = 16'b1110100111010100;
    assign mux_in_cos65 = 16'b1111111000011101;
    assign mux_in_sin65 = 16'b1110101000101011;
    assign mux_in_cos66 = 16'b1111111000001110;
    assign mux_in_sin66 = 16'b1110101010000000;
    assign mux_in_cos67 = 16'b1111110111111110;
    assign mux_in_sin67 = 16'b1110101011010100;
    assign mux_in_cos68 = 16'b1111110111101110;
    assign mux_in_sin68 = 16'b1110101100100110;
    assign mux_in_cos69 = 16'b1111110111011110;
    assign mux_in_sin69 = 16'b1110101101110111;
    assign mux_in_cos70 = 16'b1111110111001101;
    assign mux_in_sin70 = 16'b1110101111000111;
    assign mux_in_cos71 = 16'b1111110110111101;
    assign mux_in_sin71 = 16'b1110110000010110;
    assign mux_in_cos72 = 16'b1111110110101100;
    assign mux_in_sin72 = 16'b1110110001100011;
    assign mux_in_cos73 = 16'b1111110110011010;
    assign mux_in_sin73 = 16'b1110110010101111;
    assign mux_in_cos74 = 16'b1111110110001001;
    assign mux_in_sin74 = 16'b1110110011111010;
    assign mux_in_cos75 = 16'b1111110101110111;
    assign mux_in_sin75 = 16'b1110110101000100;
    assign mux_in_cos76 = 16'b1111110101100101;
    assign mux_in_sin76 = 16'b1110110110001100;
    assign mux_in_cos77 = 16'b1111110101010010;
    assign mux_in_sin77 = 16'b1110110111010100;
    assign mux_in_cos78 = 16'b1111110101000000;
    assign mux_in_sin78 = 16'b1110111000011010;
    assign mux_in_cos79 = 16'b1111110100101101;
    assign mux_in_sin79 = 16'b1110111001100000;
    assign mux_in_cos80 = 16'b1111110100011001;
    assign mux_in_sin80 = 16'b1110111010100100;
    assign mux_in_cos81 = 16'b1111110100000110;
    assign mux_in_sin81 = 16'b1110111011100111;
    assign mux_in_cos82 = 16'b1111110011110010;
    assign mux_in_sin82 = 16'b1110111100101010;
    assign mux_in_cos83 = 16'b1111110011011110;
    assign mux_in_sin83 = 16'b1110111101101011;
    assign mux_in_cos84 = 16'b1111110011001010;
    assign mux_in_sin84 = 16'b1110111110101011;
    assign mux_in_cos85 = 16'b1111110010110101;
    assign mux_in_sin85 = 16'b1110111111101011;
    assign mux_in_cos86 = 16'b1111110010100000;
    assign mux_in_sin86 = 16'b1111000000101010;
    assign mux_in_cos87 = 16'b1111110010001011;
    assign mux_in_sin87 = 16'b1111000001100111;
    assign mux_in_cos88 = 16'b1111110001110101;
    assign mux_in_sin88 = 16'b1111000010100100;
    assign mux_in_cos89 = 16'b1111110001011111;
    assign mux_in_sin89 = 16'b1111000011100000;
    assign mux_in_cos90 = 16'b1111110001001001;
    assign mux_in_sin90 = 16'b1111000100011100;
    assign mux_in_cos91 = 16'b1111110000110011;
    assign mux_in_sin91 = 16'b1111000101010110;
    assign mux_in_cos92 = 16'b1111110000011100;
    assign mux_in_sin92 = 16'b1111000110010000;
    assign mux_in_cos93 = 16'b1111110000000101;
    assign mux_in_sin93 = 16'b1111000111001001;
    assign mux_in_cos94 = 16'b1111101111101101;
    assign mux_in_sin94 = 16'b1111001000000001;
    assign mux_in_cos95 = 16'b1111101111010101;
    assign mux_in_sin95 = 16'b1111001000111000;
    assign mux_in_cos96 = 16'b1111101110111101;
    assign mux_in_sin96 = 16'b1111001001101111;
    assign mux_in_cos97 = 16'b1111101110100101;
    assign mux_in_sin97 = 16'b1111001010100101;
    assign mux_in_cos98 = 16'b1111101110001100;
    assign mux_in_sin98 = 16'b1111001011011010;
    assign mux_in_cos99 = 16'b1111101101110011;
    assign mux_in_sin99 = 16'b1111001100001110;
    assign mux_in_cos100 = 16'b1111101101011010;
    assign mux_in_sin100 = 16'b1111001101000010;
    assign mux_in_cos101 = 16'b1111101101000000;
    assign mux_in_sin101 = 16'b1111001101110101;
    assign mux_in_cos102 = 16'b1111101100100110;
    assign mux_in_sin102 = 16'b1111001110101000;
    assign mux_in_cos103 = 16'b1111101100001100;
    assign mux_in_sin103 = 16'b1111001111011010;
    assign mux_in_cos104 = 16'b1111101011110001;
    assign mux_in_sin104 = 16'b1111010000001011;
    assign mux_in_cos105 = 16'b1111101011010110;
    assign mux_in_sin105 = 16'b1111010000111011;
    assign mux_in_cos106 = 16'b1111101010111011;
    assign mux_in_sin106 = 16'b1111010001101011;
    assign mux_in_cos107 = 16'b1111101010011111;
    assign mux_in_sin107 = 16'b1111010010011011;
    assign mux_in_cos108 = 16'b1111101010000011;
    assign mux_in_sin108 = 16'b1111010011001010;
    assign mux_in_cos109 = 16'b1111101001100110;
    assign mux_in_sin109 = 16'b1111010011111000;
    assign mux_in_cos110 = 16'b1111101001001001;
    assign mux_in_sin110 = 16'b1111010100100101;
    assign mux_in_cos111 = 16'b1111101000101100;
    assign mux_in_sin111 = 16'b1111010101010010;
    assign mux_in_cos112 = 16'b1111101000001111;
    assign mux_in_sin112 = 16'b1111010101111111;
    assign mux_in_cos113 = 16'b1111100111110001;
    assign mux_in_sin113 = 16'b1111010110101011;
    assign mux_in_cos114 = 16'b1111100111010010;
    assign mux_in_sin114 = 16'b1111010111010110;
    assign mux_in_cos115 = 16'b1111100110110100;
    assign mux_in_sin115 = 16'b1111011000000001;
    assign mux_in_cos116 = 16'b1111100110010101;
    assign mux_in_sin116 = 16'b1111011000101011;
    assign mux_in_cos117 = 16'b1111100101110101;
    assign mux_in_sin117 = 16'b1111011001010101;
    assign mux_in_cos118 = 16'b1111100101010101;
    assign mux_in_sin118 = 16'b1111011001111110;
    assign mux_in_cos119 = 16'b1111100100110101;
    assign mux_in_sin119 = 16'b1111011010100111;
    assign mux_in_cos120 = 16'b1111100100010100;
    assign mux_in_sin120 = 16'b1111011011001111;
    assign mux_in_cos121 = 16'b1111100011110011;
    assign mux_in_sin121 = 16'b1111011011110111;
    assign mux_in_cos122 = 16'b1111100011010010;
    assign mux_in_sin122 = 16'b1111011100011110;
    assign mux_in_cos123 = 16'b1111100010110000;
    assign mux_in_sin123 = 16'b1111011101000101;
    assign mux_in_cos124 = 16'b1111100010001110;
    assign mux_in_sin124 = 16'b1111011101101011;
    assign mux_in_cos125 = 16'b1111100001101011;
    assign mux_in_sin125 = 16'b1111011110010001;
    assign mux_in_cos126 = 16'b1111100001001000;
    assign mux_in_sin126 = 16'b1111011110110111;
    assign mux_in_cos127 = 16'b1111100000100100;
    assign mux_in_sin127 = 16'b1111011111011100;
    assign mux_in_cos128 = 16'b1111100000000000;
    assign mux_in_sin128 = 16'b1111100000000000;
    assign mux_in_cos129 = 16'b1111011111011100;
    assign mux_in_sin129 = 16'b1111100000100100;
    assign mux_in_cos130 = 16'b1111011110110111;
    assign mux_in_sin130 = 16'b1111100001001000;
    assign mux_in_cos131 = 16'b1111011110010001;
    assign mux_in_sin131 = 16'b1111100001101011;
    assign mux_in_cos132 = 16'b1111011101101011;
    assign mux_in_sin132 = 16'b1111100010001110;
    assign mux_in_cos133 = 16'b1111011101000101;
    assign mux_in_sin133 = 16'b1111100010110000;
    assign mux_in_cos134 = 16'b1111011100011110;
    assign mux_in_sin134 = 16'b1111100011010010;
    assign mux_in_cos135 = 16'b1111011011110111;
    assign mux_in_sin135 = 16'b1111100011110011;
    assign mux_in_cos136 = 16'b1111011011001111;
    assign mux_in_sin136 = 16'b1111100100010100;
    assign mux_in_cos137 = 16'b1111011010100111;
    assign mux_in_sin137 = 16'b1111100100110101;
    assign mux_in_cos138 = 16'b1111011001111110;
    assign mux_in_sin138 = 16'b1111100101010101;
    assign mux_in_cos139 = 16'b1111011001010101;
    assign mux_in_sin139 = 16'b1111100101110101;
    assign mux_in_cos140 = 16'b1111011000101011;
    assign mux_in_sin140 = 16'b1111100110010101;
    assign mux_in_cos141 = 16'b1111011000000001;
    assign mux_in_sin141 = 16'b1111100110110100;
    assign mux_in_cos142 = 16'b1111010111010110;
    assign mux_in_sin142 = 16'b1111100111010010;
    assign mux_in_cos143 = 16'b1111010110101011;
    assign mux_in_sin143 = 16'b1111100111110001;
    assign mux_in_cos144 = 16'b1111010101111111;
    assign mux_in_sin144 = 16'b1111101000001111;
    assign mux_in_cos145 = 16'b1111010101010010;
    assign mux_in_sin145 = 16'b1111101000101100;
    assign mux_in_cos146 = 16'b1111010100100101;
    assign mux_in_sin146 = 16'b1111101001001001;
    assign mux_in_cos147 = 16'b1111010011111000;
    assign mux_in_sin147 = 16'b1111101001100110;
    assign mux_in_cos148 = 16'b1111010011001010;
    assign mux_in_sin148 = 16'b1111101010000011;
    assign mux_in_cos149 = 16'b1111010010011011;
    assign mux_in_sin149 = 16'b1111101010011111;
    assign mux_in_cos150 = 16'b1111010001101011;
    assign mux_in_sin150 = 16'b1111101010111011;
    assign mux_in_cos151 = 16'b1111010000111011;
    assign mux_in_sin151 = 16'b1111101011010110;
    assign mux_in_cos152 = 16'b1111010000001011;
    assign mux_in_sin152 = 16'b1111101011110001;
    assign mux_in_cos153 = 16'b1111001111011010;
    assign mux_in_sin153 = 16'b1111101100001100;
    assign mux_in_cos154 = 16'b1111001110101000;
    assign mux_in_sin154 = 16'b1111101100100110;
    assign mux_in_cos155 = 16'b1111001101110101;
    assign mux_in_sin155 = 16'b1111101101000000;
    assign mux_in_cos156 = 16'b1111001101000010;
    assign mux_in_sin156 = 16'b1111101101011010;
    assign mux_in_cos157 = 16'b1111001100001110;
    assign mux_in_sin157 = 16'b1111101101110011;
    assign mux_in_cos158 = 16'b1111001011011010;
    assign mux_in_sin158 = 16'b1111101110001100;
    assign mux_in_cos159 = 16'b1111001010100101;
    assign mux_in_sin159 = 16'b1111101110100101;
    assign mux_in_cos160 = 16'b1111001001101111;
    assign mux_in_sin160 = 16'b1111101110111101;
    assign mux_in_cos161 = 16'b1111001000111000;
    assign mux_in_sin161 = 16'b1111101111010101;
    assign mux_in_cos162 = 16'b1111001000000001;
    assign mux_in_sin162 = 16'b1111101111101101;
    assign mux_in_cos163 = 16'b1111000111001001;
    assign mux_in_sin163 = 16'b1111110000000101;
    assign mux_in_cos164 = 16'b1111000110010000;
    assign mux_in_sin164 = 16'b1111110000011100;
    assign mux_in_cos165 = 16'b1111000101010110;
    assign mux_in_sin165 = 16'b1111110000110011;
    assign mux_in_cos166 = 16'b1111000100011100;
    assign mux_in_sin166 = 16'b1111110001001001;
    assign mux_in_cos167 = 16'b1111000011100000;
    assign mux_in_sin167 = 16'b1111110001011111;
    assign mux_in_cos168 = 16'b1111000010100100;
    assign mux_in_sin168 = 16'b1111110001110101;
    assign mux_in_cos169 = 16'b1111000001100111;
    assign mux_in_sin169 = 16'b1111110010001011;
    assign mux_in_cos170 = 16'b1111000000101010;
    assign mux_in_sin170 = 16'b1111110010100000;
    assign mux_in_cos171 = 16'b1110111111101011;
    assign mux_in_sin171 = 16'b1111110010110101;
    assign mux_in_cos172 = 16'b1110111110101011;
    assign mux_in_sin172 = 16'b1111110011001010;
    assign mux_in_cos173 = 16'b1110111101101011;
    assign mux_in_sin173 = 16'b1111110011011110;
    assign mux_in_cos174 = 16'b1110111100101010;
    assign mux_in_sin174 = 16'b1111110011110010;
    assign mux_in_cos175 = 16'b1110111011100111;
    assign mux_in_sin175 = 16'b1111110100000110;
    assign mux_in_cos176 = 16'b1110111010100100;
    assign mux_in_sin176 = 16'b1111110100011001;
    assign mux_in_cos177 = 16'b1110111001100000;
    assign mux_in_sin177 = 16'b1111110100101101;
    assign mux_in_cos178 = 16'b1110111000011010;
    assign mux_in_sin178 = 16'b1111110101000000;
    assign mux_in_cos179 = 16'b1110110111010100;
    assign mux_in_sin179 = 16'b1111110101010010;
    assign mux_in_cos180 = 16'b1110110110001100;
    assign mux_in_sin180 = 16'b1111110101100101;
    assign mux_in_cos181 = 16'b1110110101000100;
    assign mux_in_sin181 = 16'b1111110101110111;
    assign mux_in_cos182 = 16'b1110110011111010;
    assign mux_in_sin182 = 16'b1111110110001001;
    assign mux_in_cos183 = 16'b1110110010101111;
    assign mux_in_sin183 = 16'b1111110110011010;
    assign mux_in_cos184 = 16'b1110110001100011;
    assign mux_in_sin184 = 16'b1111110110101100;
    assign mux_in_cos185 = 16'b1110110000010110;
    assign mux_in_sin185 = 16'b1111110110111101;
    assign mux_in_cos186 = 16'b1110101111000111;
    assign mux_in_sin186 = 16'b1111110111001101;
    assign mux_in_cos187 = 16'b1110101101110111;
    assign mux_in_sin187 = 16'b1111110111011110;
    assign mux_in_cos188 = 16'b1110101100100110;
    assign mux_in_sin188 = 16'b1111110111101110;
    assign mux_in_cos189 = 16'b1110101011010100;
    assign mux_in_sin189 = 16'b1111110111111110;
    assign mux_in_cos190 = 16'b1110101010000000;
    assign mux_in_sin190 = 16'b1111111000001110;
    assign mux_in_cos191 = 16'b1110101000101011;
    assign mux_in_sin191 = 16'b1111111000011101;
    assign mux_in_cos192 = 16'b1110100111010100;
    assign mux_in_sin192 = 16'b1111111000101100;
    assign mux_in_cos193 = 16'b1110100101111100;
    assign mux_in_sin193 = 16'b1111111000111011;
    assign mux_in_cos194 = 16'b1110100100100010;
    assign mux_in_sin194 = 16'b1111111001001010;
    assign mux_in_cos195 = 16'b1110100011000110;
    assign mux_in_sin195 = 16'b1111111001011000;
    assign mux_in_cos196 = 16'b1110100001101001;
    assign mux_in_sin196 = 16'b1111111001100110;
    assign mux_in_cos197 = 16'b1110100000001010;
    assign mux_in_sin197 = 16'b1111111001110100;
    assign mux_in_cos198 = 16'b1110011110101010;
    assign mux_in_sin198 = 16'b1111111010000010;
    assign mux_in_cos199 = 16'b1110011101000111;
    assign mux_in_sin199 = 16'b1111111010001111;
    assign mux_in_cos200 = 16'b1110011011100011;
    assign mux_in_sin200 = 16'b1111111010011100;
    assign mux_in_cos201 = 16'b1110011001111100;
    assign mux_in_sin201 = 16'b1111111010101001;
    assign mux_in_cos202 = 16'b1110011000010100;
    assign mux_in_sin202 = 16'b1111111010110110;
    assign mux_in_cos203 = 16'b1110010110101010;
    assign mux_in_sin203 = 16'b1111111011000010;
    assign mux_in_cos204 = 16'b1110010100111101;
    assign mux_in_sin204 = 16'b1111111011001110;
    assign mux_in_cos205 = 16'b1110010011001110;
    assign mux_in_sin205 = 16'b1111111011011010;
    assign mux_in_cos206 = 16'b1110010001011101;
    assign mux_in_sin206 = 16'b1111111011100101;
    assign mux_in_cos207 = 16'b1110001111101001;
    assign mux_in_sin207 = 16'b1111111011110001;
    assign mux_in_cos208 = 16'b1110001101110011;
    assign mux_in_sin208 = 16'b1111111011111100;
    assign mux_in_cos209 = 16'b1110001011111010;
    assign mux_in_sin209 = 16'b1111111100000111;
    assign mux_in_cos210 = 16'b1110001001111110;
    assign mux_in_sin210 = 16'b1111111100010001;
    assign mux_in_cos211 = 16'b1110001000000000;
    assign mux_in_sin211 = 16'b1111111100011100;
    assign mux_in_cos212 = 16'b1110000101111110;
    assign mux_in_sin212 = 16'b1111111100100110;
    assign mux_in_cos213 = 16'b1110000011111010;
    assign mux_in_sin213 = 16'b1111111100110000;
    assign mux_in_cos214 = 16'b1110000001110010;
    assign mux_in_sin214 = 16'b1111111100111010;
    assign mux_in_cos215 = 16'b1101111111100111;
    assign mux_in_sin215 = 16'b1111111101000011;
    assign mux_in_cos216 = 16'b1101111101011000;
    assign mux_in_sin216 = 16'b1111111101001100;
    assign mux_in_cos217 = 16'b1101111011000101;
    assign mux_in_sin217 = 16'b1111111101010101;
    assign mux_in_cos218 = 16'b1101111000101110;
    assign mux_in_sin218 = 16'b1111111101011110;
    assign mux_in_cos219 = 16'b1101110110010100;
    assign mux_in_sin219 = 16'b1111111101100110;
    assign mux_in_cos220 = 16'b1101110011110100;
    assign mux_in_sin220 = 16'b1111111101101111;
    assign mux_in_cos221 = 16'b1101110001010001;
    assign mux_in_sin221 = 16'b1111111101110111;
    assign mux_in_cos222 = 16'b1101101110101000;
    assign mux_in_sin222 = 16'b1111111101111110;
    assign mux_in_cos223 = 16'b1101101011111010;
    assign mux_in_sin223 = 16'b1111111110000110;
    assign mux_in_cos224 = 16'b1101101001000111;
    assign mux_in_sin224 = 16'b1111111110001101;
    assign mux_in_cos225 = 16'b1101100110001101;
    assign mux_in_sin225 = 16'b1111111110010100;
    assign mux_in_cos226 = 16'b1101100011001110;
    assign mux_in_sin226 = 16'b1111111110011011;
    assign mux_in_cos227 = 16'b1101100000001000;
    assign mux_in_sin227 = 16'b1111111110100010;
    assign mux_in_cos228 = 16'b1101011100111010;
    assign mux_in_sin228 = 16'b1111111110101000;
    assign mux_in_cos229 = 16'b1101011001100101;
    assign mux_in_sin229 = 16'b1111111110101111;
    assign mux_in_cos230 = 16'b1101010110001000;
    assign mux_in_sin230 = 16'b1111111110110100;
    assign mux_in_cos231 = 16'b1101010010100011;
    assign mux_in_sin231 = 16'b1111111110111010;
    assign mux_in_cos232 = 16'b1101001110110011;
    assign mux_in_sin232 = 16'b1111111111000000;
    assign mux_in_cos233 = 16'b1101001010111001;
    assign mux_in_sin233 = 16'b1111111111000101;
    assign mux_in_cos234 = 16'b1101000110110100;
    assign mux_in_sin234 = 16'b1111111111001010;
    assign mux_in_cos235 = 16'b1101000010100011;
    assign mux_in_sin235 = 16'b1111111111001111;
    assign mux_in_cos236 = 16'b1100111110000100;
    assign mux_in_sin236 = 16'b1111111111010011;
    assign mux_in_cos237 = 16'b1100111001010111;
    assign mux_in_sin237 = 16'b1111111111011000;
    assign mux_in_cos238 = 16'b1100110100011001;
    assign mux_in_sin238 = 16'b1111111111011100;
    assign mux_in_cos239 = 16'b1100101111001000;
    assign mux_in_sin239 = 16'b1111111111100000;
    assign mux_in_cos240 = 16'b1100101001100011;
    assign mux_in_sin240 = 16'b1111111111100011;
    assign mux_in_cos241 = 16'b1100100011100111;
    assign mux_in_sin241 = 16'b1111111111100111;
    assign mux_in_cos242 = 16'b1100011101010000;
    assign mux_in_sin242 = 16'b1111111111101010;
    assign mux_in_cos243 = 16'b1100010110011011;
    assign mux_in_sin243 = 16'b1111111111101101;
    assign mux_in_cos244 = 16'b1100001111000011;
    assign mux_in_sin244 = 16'b1111111111110000;
    assign mux_in_cos245 = 16'b1100000111000010;
    assign mux_in_sin245 = 16'b1111111111110011;
    assign mux_in_cos246 = 16'b1011111110001111;
    assign mux_in_sin246 = 16'b1111111111110101;
    assign mux_in_cos247 = 16'b1011110100100010;
    assign mux_in_sin247 = 16'b1111111111110111;
    assign mux_in_cos248 = 16'b1011101001101010;
    assign mux_in_sin248 = 16'b1111111111111001;
    assign mux_in_cos249 = 16'b1011011101010110;
    assign mux_in_sin249 = 16'b1111111111111011;
    assign mux_in_cos250 = 16'b1011001111000111;
    assign mux_in_sin250 = 16'b1111111111111100;
    assign mux_in_cos251 = 16'b1010111110010010;
    assign mux_in_sin251 = 16'b1111111111111101;
    assign mux_in_cos252 = 16'b1010101001101100;
    assign mux_in_sin252 = 16'b1111111111111110;
    assign mux_in_cos253 = 16'b1010001111001000;
    assign mux_in_sin253 = 16'b1111111111111111;
    assign mux_in_cos254 = 16'b1001101001101100;
    assign mux_in_sin254 = 16'b0000000000000000;
    assign mux_in_cos255 = 16'b1000101001101100;
    assign mux_in_sin255 = 16'b0000000000000000;
    assign mux_in_cos256 = 16'b0000000000000000;
    assign mux_in_sin256 = 16'b0000000000000000;

    always @ (*)
    begin
        case(x_in1)
        9'b000000000 : logsin1 = mux_in_sin0;
        9'b000000001 : logsin1 = mux_in_sin1;
        9'b000000010 : logsin1 = mux_in_sin2;
        9'b000000011 : logsin1 = mux_in_sin3;
        9'b000000100 : logsin1 = mux_in_sin4;
        9'b000000101 : logsin1 = mux_in_sin5;
        9'b000000110 : logsin1 = mux_in_sin6;
        9'b000000111 : logsin1 = mux_in_sin7;
        9'b000001000 : logsin1 = mux_in_sin8;
        9'b000001001 : logsin1 = mux_in_sin9;
        9'b000001010 : logsin1 = mux_in_sin10;
        9'b000001011 : logsin1 = mux_in_sin11;
        9'b000001100 : logsin1 = mux_in_sin12;
        9'b000001101 : logsin1 = mux_in_sin13;
        9'b000001110 : logsin1 = mux_in_sin14;
        9'b000001111 : logsin1 = mux_in_sin15;
        9'b000010000 : logsin1 = mux_in_sin16;
        9'b000010001 : logsin1 = mux_in_sin17;
        9'b000010010 : logsin1 = mux_in_sin18;
        9'b000010011 : logsin1 = mux_in_sin19;
        9'b000010100 : logsin1 = mux_in_sin20;
        9'b000010101 : logsin1 = mux_in_sin21;
        9'b000010110 : logsin1 = mux_in_sin22;
        9'b000010111 : logsin1 = mux_in_sin23;
        9'b000011000 : logsin1 = mux_in_sin24;
        9'b000011001 : logsin1 = mux_in_sin25;
        9'b000011010 : logsin1 = mux_in_sin26;
        9'b000011011 : logsin1 = mux_in_sin27;
        9'b000011100 : logsin1 = mux_in_sin28;
        9'b000011101 : logsin1 = mux_in_sin29;
        9'b000011110 : logsin1 = mux_in_sin30;
        9'b000011111 : logsin1 = mux_in_sin31;
        9'b000100000 : logsin1 = mux_in_sin32;
        9'b000100001 : logsin1 = mux_in_sin33;
        9'b000100010 : logsin1 = mux_in_sin34;
        9'b000100011 : logsin1 = mux_in_sin35;
        9'b000100100 : logsin1 = mux_in_sin36;
        9'b000100101 : logsin1 = mux_in_sin37;
        9'b000100110 : logsin1 = mux_in_sin38;
        9'b000100111 : logsin1 = mux_in_sin39;
        9'b000101000 : logsin1 = mux_in_sin40;
        9'b000101001 : logsin1 = mux_in_sin41;
        9'b000101010 : logsin1 = mux_in_sin42;
        9'b000101011 : logsin1 = mux_in_sin43;
        9'b000101100 : logsin1 = mux_in_sin44;
        9'b000101101 : logsin1 = mux_in_sin45;
        9'b000101110 : logsin1 = mux_in_sin46;
        9'b000101111 : logsin1 = mux_in_sin47;
        9'b000110000 : logsin1 = mux_in_sin48;
        9'b000110001 : logsin1 = mux_in_sin49;
        9'b000110010 : logsin1 = mux_in_sin50;
        9'b000110011 : logsin1 = mux_in_sin51;
        9'b000110100 : logsin1 = mux_in_sin52;
        9'b000110101 : logsin1 = mux_in_sin53;
        9'b000110110 : logsin1 = mux_in_sin54;
        9'b000110111 : logsin1 = mux_in_sin55;
        9'b000111000 : logsin1 = mux_in_sin56;
        9'b000111001 : logsin1 = mux_in_sin57;
        9'b000111010 : logsin1 = mux_in_sin58;
        9'b000111011 : logsin1 = mux_in_sin59;
        9'b000111100 : logsin1 = mux_in_sin60;
        9'b000111101 : logsin1 = mux_in_sin61;
        9'b000111110 : logsin1 = mux_in_sin62;
        9'b000111111 : logsin1 = mux_in_sin63;
        9'b001000000 : logsin1 = mux_in_sin64;
        9'b001000001 : logsin1 = mux_in_sin65;
        9'b001000010 : logsin1 = mux_in_sin66;
        9'b001000011 : logsin1 = mux_in_sin67;
        9'b001000100 : logsin1 = mux_in_sin68;
        9'b001000101 : logsin1 = mux_in_sin69;
        9'b001000110 : logsin1 = mux_in_sin70;
        9'b001000111 : logsin1 = mux_in_sin71;
        9'b001001000 : logsin1 = mux_in_sin72;
        9'b001001001 : logsin1 = mux_in_sin73;
        9'b001001010 : logsin1 = mux_in_sin74;
        9'b001001011 : logsin1 = mux_in_sin75;
        9'b001001100 : logsin1 = mux_in_sin76;
        9'b001001101 : logsin1 = mux_in_sin77;
        9'b001001110 : logsin1 = mux_in_sin78;
        9'b001001111 : logsin1 = mux_in_sin79;
        9'b001010000 : logsin1 = mux_in_sin80;
        9'b001010001 : logsin1 = mux_in_sin81;
        9'b001010010 : logsin1 = mux_in_sin82;
        9'b001010011 : logsin1 = mux_in_sin83;
        9'b001010100 : logsin1 = mux_in_sin84;
        9'b001010101 : logsin1 = mux_in_sin85;
        9'b001010110 : logsin1 = mux_in_sin86;
        9'b001010111 : logsin1 = mux_in_sin87;
        9'b001011000 : logsin1 = mux_in_sin88;
        9'b001011001 : logsin1 = mux_in_sin89;
        9'b001011010 : logsin1 = mux_in_sin90;
        9'b001011011 : logsin1 = mux_in_sin91;
        9'b001011100 : logsin1 = mux_in_sin92;
        9'b001011101 : logsin1 = mux_in_sin93;
        9'b001011110 : logsin1 = mux_in_sin94;
        9'b001011111 : logsin1 = mux_in_sin95;
        9'b001100000 : logsin1 = mux_in_sin96;
        9'b001100001 : logsin1 = mux_in_sin97;
        9'b001100010 : logsin1 = mux_in_sin98;
        9'b001100011 : logsin1 = mux_in_sin99;
        9'b001100100 : logsin1 = mux_in_sin100;
        9'b001100101 : logsin1 = mux_in_sin101;
        9'b001100110 : logsin1 = mux_in_sin102;
        9'b001100111 : logsin1 = mux_in_sin103;
        9'b001101000 : logsin1 = mux_in_sin104;
        9'b001101001 : logsin1 = mux_in_sin105;
        9'b001101010 : logsin1 = mux_in_sin106;
        9'b001101011 : logsin1 = mux_in_sin107;
        9'b001101100 : logsin1 = mux_in_sin108;
        9'b001101101 : logsin1 = mux_in_sin109;
        9'b001101110 : logsin1 = mux_in_sin110;
        9'b001101111 : logsin1 = mux_in_sin111;
        9'b001110000 : logsin1 = mux_in_sin112;
        9'b001110001 : logsin1 = mux_in_sin113;
        9'b001110010 : logsin1 = mux_in_sin114;
        9'b001110011 : logsin1 = mux_in_sin115;
        9'b001110100 : logsin1 = mux_in_sin116;
        9'b001110101 : logsin1 = mux_in_sin117;
        9'b001110110 : logsin1 = mux_in_sin118;
        9'b001110111 : logsin1 = mux_in_sin119;
        9'b001111000 : logsin1 = mux_in_sin120;
        9'b001111001 : logsin1 = mux_in_sin121;
        9'b001111010 : logsin1 = mux_in_sin122;
        9'b001111011 : logsin1 = mux_in_sin123;
        9'b001111100 : logsin1 = mux_in_sin124;
        9'b001111101 : logsin1 = mux_in_sin125;
        9'b001111110 : logsin1 = mux_in_sin126;
        9'b001111111 : logsin1 = mux_in_sin127;
        9'b010000000 : logsin1 = mux_in_sin128;
        9'b010000001 : logsin1 = mux_in_sin129;
        9'b010000010 : logsin1 = mux_in_sin130;
        9'b010000011 : logsin1 = mux_in_sin131;
        9'b010000100 : logsin1 = mux_in_sin132;
        9'b010000101 : logsin1 = mux_in_sin133;
        9'b010000110 : logsin1 = mux_in_sin134;
        9'b010000111 : logsin1 = mux_in_sin135;
        9'b010001000 : logsin1 = mux_in_sin136;
        9'b010001001 : logsin1 = mux_in_sin137;
        9'b010001010 : logsin1 = mux_in_sin138;
        9'b010001011 : logsin1 = mux_in_sin139;
        9'b010001100 : logsin1 = mux_in_sin140;
        9'b010001101 : logsin1 = mux_in_sin141;
        9'b010001110 : logsin1 = mux_in_sin142;
        9'b010001111 : logsin1 = mux_in_sin143;
        9'b010010000 : logsin1 = mux_in_sin144;
        9'b010010001 : logsin1 = mux_in_sin145;
        9'b010010010 : logsin1 = mux_in_sin146;
        9'b010010011 : logsin1 = mux_in_sin147;
        9'b010010100 : logsin1 = mux_in_sin148;
        9'b010010101 : logsin1 = mux_in_sin149;
        9'b010010110 : logsin1 = mux_in_sin150;
        9'b010010111 : logsin1 = mux_in_sin151;
        9'b010011000 : logsin1 = mux_in_sin152;
        9'b010011001 : logsin1 = mux_in_sin153;
        9'b010011010 : logsin1 = mux_in_sin154;
        9'b010011011 : logsin1 = mux_in_sin155;
        9'b010011100 : logsin1 = mux_in_sin156;
        9'b010011101 : logsin1 = mux_in_sin157;
        9'b010011110 : logsin1 = mux_in_sin158;
        9'b010011111 : logsin1 = mux_in_sin159;
        9'b010100000 : logsin1 = mux_in_sin160;
        9'b010100001 : logsin1 = mux_in_sin161;
        9'b010100010 : logsin1 = mux_in_sin162;
        9'b010100011 : logsin1 = mux_in_sin163;
        9'b010100100 : logsin1 = mux_in_sin164;
        9'b010100101 : logsin1 = mux_in_sin165;
        9'b010100110 : logsin1 = mux_in_sin166;
        9'b010100111 : logsin1 = mux_in_sin167;
        9'b010101000 : logsin1 = mux_in_sin168;
        9'b010101001 : logsin1 = mux_in_sin169;
        9'b010101010 : logsin1 = mux_in_sin170;
        9'b010101011 : logsin1 = mux_in_sin171;
        9'b010101100 : logsin1 = mux_in_sin172;
        9'b010101101 : logsin1 = mux_in_sin173;
        9'b010101110 : logsin1 = mux_in_sin174;
        9'b010101111 : logsin1 = mux_in_sin175;
        9'b010110000 : logsin1 = mux_in_sin176;
        9'b010110001 : logsin1 = mux_in_sin177;
        9'b010110010 : logsin1 = mux_in_sin178;
        9'b010110011 : logsin1 = mux_in_sin179;
        9'b010110100 : logsin1 = mux_in_sin180;
        9'b010110101 : logsin1 = mux_in_sin181;
        9'b010110110 : logsin1 = mux_in_sin182;
        9'b010110111 : logsin1 = mux_in_sin183;
        9'b010111000 : logsin1 = mux_in_sin184;
        9'b010111001 : logsin1 = mux_in_sin185;
        9'b010111010 : logsin1 = mux_in_sin186;
        9'b010111011 : logsin1 = mux_in_sin187;
        9'b010111100 : logsin1 = mux_in_sin188;
        9'b010111101 : logsin1 = mux_in_sin189;
        9'b010111110 : logsin1 = mux_in_sin190;
        9'b010111111 : logsin1 = mux_in_sin191;
        9'b011000000 : logsin1 = mux_in_sin192;
        9'b011000001 : logsin1 = mux_in_sin193;
        9'b011000010 : logsin1 = mux_in_sin194;
        9'b011000011 : logsin1 = mux_in_sin195;
        9'b011000100 : logsin1 = mux_in_sin196;
        9'b011000101 : logsin1 = mux_in_sin197;
        9'b011000110 : logsin1 = mux_in_sin198;
        9'b011000111 : logsin1 = mux_in_sin199;
        9'b011001000 : logsin1 = mux_in_sin200;
        9'b011001001 : logsin1 = mux_in_sin201;
        9'b011001010 : logsin1 = mux_in_sin202;
        9'b011001011 : logsin1 = mux_in_sin203;
        9'b011001100 : logsin1 = mux_in_sin204;
        9'b011001101 : logsin1 = mux_in_sin205;
        9'b011001110 : logsin1 = mux_in_sin206;
        9'b011001111 : logsin1 = mux_in_sin207;
        9'b011010000 : logsin1 = mux_in_sin208;
        9'b011010001 : logsin1 = mux_in_sin209;
        9'b011010010 : logsin1 = mux_in_sin210;
        9'b011010011 : logsin1 = mux_in_sin211;
        9'b011010100 : logsin1 = mux_in_sin212;
        9'b011010101 : logsin1 = mux_in_sin213;
        9'b011010110 : logsin1 = mux_in_sin214;
        9'b011010111 : logsin1 = mux_in_sin215;
        9'b011011000 : logsin1 = mux_in_sin216;
        9'b011011001 : logsin1 = mux_in_sin217;
        9'b011011010 : logsin1 = mux_in_sin218;
        9'b011011011 : logsin1 = mux_in_sin219;
        9'b011011100 : logsin1 = mux_in_sin220;
        9'b011011101 : logsin1 = mux_in_sin221;
        9'b011011110 : logsin1 = mux_in_sin222;
        9'b011011111 : logsin1 = mux_in_sin223;
        9'b011100000 : logsin1 = mux_in_sin224;
        9'b011100001 : logsin1 = mux_in_sin225;
        9'b011100010 : logsin1 = mux_in_sin226;
        9'b011100011 : logsin1 = mux_in_sin227;
        9'b011100100 : logsin1 = mux_in_sin228;
        9'b011100101 : logsin1 = mux_in_sin229;
        9'b011100110 : logsin1 = mux_in_sin230;
        9'b011100111 : logsin1 = mux_in_sin231;
        9'b011101000 : logsin1 = mux_in_sin232;
        9'b011101001 : logsin1 = mux_in_sin233;
        9'b011101010 : logsin1 = mux_in_sin234;
        9'b011101011 : logsin1 = mux_in_sin235;
        9'b011101100 : logsin1 = mux_in_sin236;
        9'b011101101 : logsin1 = mux_in_sin237;
        9'b011101110 : logsin1 = mux_in_sin238;
        9'b011101111 : logsin1 = mux_in_sin239;
        9'b011110000 : logsin1 = mux_in_sin240;
        9'b011110001 : logsin1 = mux_in_sin241;
        9'b011110010 : logsin1 = mux_in_sin242;
        9'b011110011 : logsin1 = mux_in_sin243;
        9'b011110100 : logsin1 = mux_in_sin244;
        9'b011110101 : logsin1 = mux_in_sin245;
        9'b011110110 : logsin1 = mux_in_sin246;
        9'b011110111 : logsin1 = mux_in_sin247;
        9'b011111000 : logsin1 = mux_in_sin248;
        9'b011111001 : logsin1 = mux_in_sin249;
        9'b011111010 : logsin1 = mux_in_sin250;
        9'b011111011 : logsin1 = mux_in_sin251;
        9'b011111100 : logsin1 = mux_in_sin252;
        9'b011111101 : logsin1 = mux_in_sin253;
        9'b011111110 : logsin1 = mux_in_sin254;
        9'b011111111 : logsin1 = mux_in_sin255;
        9'b100000000 : logsin1 = mux_in_sin256;
        default: logsin1 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in2)
        9'b000000000 : logsin2 = mux_in_sin0;
        9'b000000001 : logsin2 = mux_in_sin1;
        9'b000000010 : logsin2 = mux_in_sin2;
        9'b000000011 : logsin2 = mux_in_sin3;
        9'b000000100 : logsin2 = mux_in_sin4;
        9'b000000101 : logsin2 = mux_in_sin5;
        9'b000000110 : logsin2 = mux_in_sin6;
        9'b000000111 : logsin2 = mux_in_sin7;
        9'b000001000 : logsin2 = mux_in_sin8;
        9'b000001001 : logsin2 = mux_in_sin9;
        9'b000001010 : logsin2 = mux_in_sin10;
        9'b000001011 : logsin2 = mux_in_sin11;
        9'b000001100 : logsin2 = mux_in_sin12;
        9'b000001101 : logsin2 = mux_in_sin13;
        9'b000001110 : logsin2 = mux_in_sin14;
        9'b000001111 : logsin2 = mux_in_sin15;
        9'b000010000 : logsin2 = mux_in_sin16;
        9'b000010001 : logsin2 = mux_in_sin17;
        9'b000010010 : logsin2 = mux_in_sin18;
        9'b000010011 : logsin2 = mux_in_sin19;
        9'b000010100 : logsin2 = mux_in_sin20;
        9'b000010101 : logsin2 = mux_in_sin21;
        9'b000010110 : logsin2 = mux_in_sin22;
        9'b000010111 : logsin2 = mux_in_sin23;
        9'b000011000 : logsin2 = mux_in_sin24;
        9'b000011001 : logsin2 = mux_in_sin25;
        9'b000011010 : logsin2 = mux_in_sin26;
        9'b000011011 : logsin2 = mux_in_sin27;
        9'b000011100 : logsin2 = mux_in_sin28;
        9'b000011101 : logsin2 = mux_in_sin29;
        9'b000011110 : logsin2 = mux_in_sin30;
        9'b000011111 : logsin2 = mux_in_sin31;
        9'b000100000 : logsin2 = mux_in_sin32;
        9'b000100001 : logsin2 = mux_in_sin33;
        9'b000100010 : logsin2 = mux_in_sin34;
        9'b000100011 : logsin2 = mux_in_sin35;
        9'b000100100 : logsin2 = mux_in_sin36;
        9'b000100101 : logsin2 = mux_in_sin37;
        9'b000100110 : logsin2 = mux_in_sin38;
        9'b000100111 : logsin2 = mux_in_sin39;
        9'b000101000 : logsin2 = mux_in_sin40;
        9'b000101001 : logsin2 = mux_in_sin41;
        9'b000101010 : logsin2 = mux_in_sin42;
        9'b000101011 : logsin2 = mux_in_sin43;
        9'b000101100 : logsin2 = mux_in_sin44;
        9'b000101101 : logsin2 = mux_in_sin45;
        9'b000101110 : logsin2 = mux_in_sin46;
        9'b000101111 : logsin2 = mux_in_sin47;
        9'b000110000 : logsin2 = mux_in_sin48;
        9'b000110001 : logsin2 = mux_in_sin49;
        9'b000110010 : logsin2 = mux_in_sin50;
        9'b000110011 : logsin2 = mux_in_sin51;
        9'b000110100 : logsin2 = mux_in_sin52;
        9'b000110101 : logsin2 = mux_in_sin53;
        9'b000110110 : logsin2 = mux_in_sin54;
        9'b000110111 : logsin2 = mux_in_sin55;
        9'b000111000 : logsin2 = mux_in_sin56;
        9'b000111001 : logsin2 = mux_in_sin57;
        9'b000111010 : logsin2 = mux_in_sin58;
        9'b000111011 : logsin2 = mux_in_sin59;
        9'b000111100 : logsin2 = mux_in_sin60;
        9'b000111101 : logsin2 = mux_in_sin61;
        9'b000111110 : logsin2 = mux_in_sin62;
        9'b000111111 : logsin2 = mux_in_sin63;
        9'b001000000 : logsin2 = mux_in_sin64;
        9'b001000001 : logsin2 = mux_in_sin65;
        9'b001000010 : logsin2 = mux_in_sin66;
        9'b001000011 : logsin2 = mux_in_sin67;
        9'b001000100 : logsin2 = mux_in_sin68;
        9'b001000101 : logsin2 = mux_in_sin69;
        9'b001000110 : logsin2 = mux_in_sin70;
        9'b001000111 : logsin2 = mux_in_sin71;
        9'b001001000 : logsin2 = mux_in_sin72;
        9'b001001001 : logsin2 = mux_in_sin73;
        9'b001001010 : logsin2 = mux_in_sin74;
        9'b001001011 : logsin2 = mux_in_sin75;
        9'b001001100 : logsin2 = mux_in_sin76;
        9'b001001101 : logsin2 = mux_in_sin77;
        9'b001001110 : logsin2 = mux_in_sin78;
        9'b001001111 : logsin2 = mux_in_sin79;
        9'b001010000 : logsin2 = mux_in_sin80;
        9'b001010001 : logsin2 = mux_in_sin81;
        9'b001010010 : logsin2 = mux_in_sin82;
        9'b001010011 : logsin2 = mux_in_sin83;
        9'b001010100 : logsin2 = mux_in_sin84;
        9'b001010101 : logsin2 = mux_in_sin85;
        9'b001010110 : logsin2 = mux_in_sin86;
        9'b001010111 : logsin2 = mux_in_sin87;
        9'b001011000 : logsin2 = mux_in_sin88;
        9'b001011001 : logsin2 = mux_in_sin89;
        9'b001011010 : logsin2 = mux_in_sin90;
        9'b001011011 : logsin2 = mux_in_sin91;
        9'b001011100 : logsin2 = mux_in_sin92;
        9'b001011101 : logsin2 = mux_in_sin93;
        9'b001011110 : logsin2 = mux_in_sin94;
        9'b001011111 : logsin2 = mux_in_sin95;
        9'b001100000 : logsin2 = mux_in_sin96;
        9'b001100001 : logsin2 = mux_in_sin97;
        9'b001100010 : logsin2 = mux_in_sin98;
        9'b001100011 : logsin2 = mux_in_sin99;
        9'b001100100 : logsin2 = mux_in_sin100;
        9'b001100101 : logsin2 = mux_in_sin101;
        9'b001100110 : logsin2 = mux_in_sin102;
        9'b001100111 : logsin2 = mux_in_sin103;
        9'b001101000 : logsin2 = mux_in_sin104;
        9'b001101001 : logsin2 = mux_in_sin105;
        9'b001101010 : logsin2 = mux_in_sin106;
        9'b001101011 : logsin2 = mux_in_sin107;
        9'b001101100 : logsin2 = mux_in_sin108;
        9'b001101101 : logsin2 = mux_in_sin109;
        9'b001101110 : logsin2 = mux_in_sin110;
        9'b001101111 : logsin2 = mux_in_sin111;
        9'b001110000 : logsin2 = mux_in_sin112;
        9'b001110001 : logsin2 = mux_in_sin113;
        9'b001110010 : logsin2 = mux_in_sin114;
        9'b001110011 : logsin2 = mux_in_sin115;
        9'b001110100 : logsin2 = mux_in_sin116;
        9'b001110101 : logsin2 = mux_in_sin117;
        9'b001110110 : logsin2 = mux_in_sin118;
        9'b001110111 : logsin2 = mux_in_sin119;
        9'b001111000 : logsin2 = mux_in_sin120;
        9'b001111001 : logsin2 = mux_in_sin121;
        9'b001111010 : logsin2 = mux_in_sin122;
        9'b001111011 : logsin2 = mux_in_sin123;
        9'b001111100 : logsin2 = mux_in_sin124;
        9'b001111101 : logsin2 = mux_in_sin125;
        9'b001111110 : logsin2 = mux_in_sin126;
        9'b001111111 : logsin2 = mux_in_sin127;
        9'b010000000 : logsin2 = mux_in_sin128;
        9'b010000001 : logsin2 = mux_in_sin129;
        9'b010000010 : logsin2 = mux_in_sin130;
        9'b010000011 : logsin2 = mux_in_sin131;
        9'b010000100 : logsin2 = mux_in_sin132;
        9'b010000101 : logsin2 = mux_in_sin133;
        9'b010000110 : logsin2 = mux_in_sin134;
        9'b010000111 : logsin2 = mux_in_sin135;
        9'b010001000 : logsin2 = mux_in_sin136;
        9'b010001001 : logsin2 = mux_in_sin137;
        9'b010001010 : logsin2 = mux_in_sin138;
        9'b010001011 : logsin2 = mux_in_sin139;
        9'b010001100 : logsin2 = mux_in_sin140;
        9'b010001101 : logsin2 = mux_in_sin141;
        9'b010001110 : logsin2 = mux_in_sin142;
        9'b010001111 : logsin2 = mux_in_sin143;
        9'b010010000 : logsin2 = mux_in_sin144;
        9'b010010001 : logsin2 = mux_in_sin145;
        9'b010010010 : logsin2 = mux_in_sin146;
        9'b010010011 : logsin2 = mux_in_sin147;
        9'b010010100 : logsin2 = mux_in_sin148;
        9'b010010101 : logsin2 = mux_in_sin149;
        9'b010010110 : logsin2 = mux_in_sin150;
        9'b010010111 : logsin2 = mux_in_sin151;
        9'b010011000 : logsin2 = mux_in_sin152;
        9'b010011001 : logsin2 = mux_in_sin153;
        9'b010011010 : logsin2 = mux_in_sin154;
        9'b010011011 : logsin2 = mux_in_sin155;
        9'b010011100 : logsin2 = mux_in_sin156;
        9'b010011101 : logsin2 = mux_in_sin157;
        9'b010011110 : logsin2 = mux_in_sin158;
        9'b010011111 : logsin2 = mux_in_sin159;
        9'b010100000 : logsin2 = mux_in_sin160;
        9'b010100001 : logsin2 = mux_in_sin161;
        9'b010100010 : logsin2 = mux_in_sin162;
        9'b010100011 : logsin2 = mux_in_sin163;
        9'b010100100 : logsin2 = mux_in_sin164;
        9'b010100101 : logsin2 = mux_in_sin165;
        9'b010100110 : logsin2 = mux_in_sin166;
        9'b010100111 : logsin2 = mux_in_sin167;
        9'b010101000 : logsin2 = mux_in_sin168;
        9'b010101001 : logsin2 = mux_in_sin169;
        9'b010101010 : logsin2 = mux_in_sin170;
        9'b010101011 : logsin2 = mux_in_sin171;
        9'b010101100 : logsin2 = mux_in_sin172;
        9'b010101101 : logsin2 = mux_in_sin173;
        9'b010101110 : logsin2 = mux_in_sin174;
        9'b010101111 : logsin2 = mux_in_sin175;
        9'b010110000 : logsin2 = mux_in_sin176;
        9'b010110001 : logsin2 = mux_in_sin177;
        9'b010110010 : logsin2 = mux_in_sin178;
        9'b010110011 : logsin2 = mux_in_sin179;
        9'b010110100 : logsin2 = mux_in_sin180;
        9'b010110101 : logsin2 = mux_in_sin181;
        9'b010110110 : logsin2 = mux_in_sin182;
        9'b010110111 : logsin2 = mux_in_sin183;
        9'b010111000 : logsin2 = mux_in_sin184;
        9'b010111001 : logsin2 = mux_in_sin185;
        9'b010111010 : logsin2 = mux_in_sin186;
        9'b010111011 : logsin2 = mux_in_sin187;
        9'b010111100 : logsin2 = mux_in_sin188;
        9'b010111101 : logsin2 = mux_in_sin189;
        9'b010111110 : logsin2 = mux_in_sin190;
        9'b010111111 : logsin2 = mux_in_sin191;
        9'b011000000 : logsin2 = mux_in_sin192;
        9'b011000001 : logsin2 = mux_in_sin193;
        9'b011000010 : logsin2 = mux_in_sin194;
        9'b011000011 : logsin2 = mux_in_sin195;
        9'b011000100 : logsin2 = mux_in_sin196;
        9'b011000101 : logsin2 = mux_in_sin197;
        9'b011000110 : logsin2 = mux_in_sin198;
        9'b011000111 : logsin2 = mux_in_sin199;
        9'b011001000 : logsin2 = mux_in_sin200;
        9'b011001001 : logsin2 = mux_in_sin201;
        9'b011001010 : logsin2 = mux_in_sin202;
        9'b011001011 : logsin2 = mux_in_sin203;
        9'b011001100 : logsin2 = mux_in_sin204;
        9'b011001101 : logsin2 = mux_in_sin205;
        9'b011001110 : logsin2 = mux_in_sin206;
        9'b011001111 : logsin2 = mux_in_sin207;
        9'b011010000 : logsin2 = mux_in_sin208;
        9'b011010001 : logsin2 = mux_in_sin209;
        9'b011010010 : logsin2 = mux_in_sin210;
        9'b011010011 : logsin2 = mux_in_sin211;
        9'b011010100 : logsin2 = mux_in_sin212;
        9'b011010101 : logsin2 = mux_in_sin213;
        9'b011010110 : logsin2 = mux_in_sin214;
        9'b011010111 : logsin2 = mux_in_sin215;
        9'b011011000 : logsin2 = mux_in_sin216;
        9'b011011001 : logsin2 = mux_in_sin217;
        9'b011011010 : logsin2 = mux_in_sin218;
        9'b011011011 : logsin2 = mux_in_sin219;
        9'b011011100 : logsin2 = mux_in_sin220;
        9'b011011101 : logsin2 = mux_in_sin221;
        9'b011011110 : logsin2 = mux_in_sin222;
        9'b011011111 : logsin2 = mux_in_sin223;
        9'b011100000 : logsin2 = mux_in_sin224;
        9'b011100001 : logsin2 = mux_in_sin225;
        9'b011100010 : logsin2 = mux_in_sin226;
        9'b011100011 : logsin2 = mux_in_sin227;
        9'b011100100 : logsin2 = mux_in_sin228;
        9'b011100101 : logsin2 = mux_in_sin229;
        9'b011100110 : logsin2 = mux_in_sin230;
        9'b011100111 : logsin2 = mux_in_sin231;
        9'b011101000 : logsin2 = mux_in_sin232;
        9'b011101001 : logsin2 = mux_in_sin233;
        9'b011101010 : logsin2 = mux_in_sin234;
        9'b011101011 : logsin2 = mux_in_sin235;
        9'b011101100 : logsin2 = mux_in_sin236;
        9'b011101101 : logsin2 = mux_in_sin237;
        9'b011101110 : logsin2 = mux_in_sin238;
        9'b011101111 : logsin2 = mux_in_sin239;
        9'b011110000 : logsin2 = mux_in_sin240;
        9'b011110001 : logsin2 = mux_in_sin241;
        9'b011110010 : logsin2 = mux_in_sin242;
        9'b011110011 : logsin2 = mux_in_sin243;
        9'b011110100 : logsin2 = mux_in_sin244;
        9'b011110101 : logsin2 = mux_in_sin245;
        9'b011110110 : logsin2 = mux_in_sin246;
        9'b011110111 : logsin2 = mux_in_sin247;
        9'b011111000 : logsin2 = mux_in_sin248;
        9'b011111001 : logsin2 = mux_in_sin249;
        9'b011111010 : logsin2 = mux_in_sin250;
        9'b011111011 : logsin2 = mux_in_sin251;
        9'b011111100 : logsin2 = mux_in_sin252;
        9'b011111101 : logsin2 = mux_in_sin253;
        9'b011111110 : logsin2 = mux_in_sin254;
        9'b011111111 : logsin2 = mux_in_sin255;
        9'b100000000 : logsin2 = mux_in_sin256;
        default: logsin2 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in3)
        9'b000000000 : logsin3 = mux_in_sin0;
        9'b000000001 : logsin3 = mux_in_sin1;
        9'b000000010 : logsin3 = mux_in_sin2;
        9'b000000011 : logsin3 = mux_in_sin3;
        9'b000000100 : logsin3 = mux_in_sin4;
        9'b000000101 : logsin3 = mux_in_sin5;
        9'b000000110 : logsin3 = mux_in_sin6;
        9'b000000111 : logsin3 = mux_in_sin7;
        9'b000001000 : logsin3 = mux_in_sin8;
        9'b000001001 : logsin3 = mux_in_sin9;
        9'b000001010 : logsin3 = mux_in_sin10;
        9'b000001011 : logsin3 = mux_in_sin11;
        9'b000001100 : logsin3 = mux_in_sin12;
        9'b000001101 : logsin3 = mux_in_sin13;
        9'b000001110 : logsin3 = mux_in_sin14;
        9'b000001111 : logsin3 = mux_in_sin15;
        9'b000010000 : logsin3 = mux_in_sin16;
        9'b000010001 : logsin3 = mux_in_sin17;
        9'b000010010 : logsin3 = mux_in_sin18;
        9'b000010011 : logsin3 = mux_in_sin19;
        9'b000010100 : logsin3 = mux_in_sin20;
        9'b000010101 : logsin3 = mux_in_sin21;
        9'b000010110 : logsin3 = mux_in_sin22;
        9'b000010111 : logsin3 = mux_in_sin23;
        9'b000011000 : logsin3 = mux_in_sin24;
        9'b000011001 : logsin3 = mux_in_sin25;
        9'b000011010 : logsin3 = mux_in_sin26;
        9'b000011011 : logsin3 = mux_in_sin27;
        9'b000011100 : logsin3 = mux_in_sin28;
        9'b000011101 : logsin3 = mux_in_sin29;
        9'b000011110 : logsin3 = mux_in_sin30;
        9'b000011111 : logsin3 = mux_in_sin31;
        9'b000100000 : logsin3 = mux_in_sin32;
        9'b000100001 : logsin3 = mux_in_sin33;
        9'b000100010 : logsin3 = mux_in_sin34;
        9'b000100011 : logsin3 = mux_in_sin35;
        9'b000100100 : logsin3 = mux_in_sin36;
        9'b000100101 : logsin3 = mux_in_sin37;
        9'b000100110 : logsin3 = mux_in_sin38;
        9'b000100111 : logsin3 = mux_in_sin39;
        9'b000101000 : logsin3 = mux_in_sin40;
        9'b000101001 : logsin3 = mux_in_sin41;
        9'b000101010 : logsin3 = mux_in_sin42;
        9'b000101011 : logsin3 = mux_in_sin43;
        9'b000101100 : logsin3 = mux_in_sin44;
        9'b000101101 : logsin3 = mux_in_sin45;
        9'b000101110 : logsin3 = mux_in_sin46;
        9'b000101111 : logsin3 = mux_in_sin47;
        9'b000110000 : logsin3 = mux_in_sin48;
        9'b000110001 : logsin3 = mux_in_sin49;
        9'b000110010 : logsin3 = mux_in_sin50;
        9'b000110011 : logsin3 = mux_in_sin51;
        9'b000110100 : logsin3 = mux_in_sin52;
        9'b000110101 : logsin3 = mux_in_sin53;
        9'b000110110 : logsin3 = mux_in_sin54;
        9'b000110111 : logsin3 = mux_in_sin55;
        9'b000111000 : logsin3 = mux_in_sin56;
        9'b000111001 : logsin3 = mux_in_sin57;
        9'b000111010 : logsin3 = mux_in_sin58;
        9'b000111011 : logsin3 = mux_in_sin59;
        9'b000111100 : logsin3 = mux_in_sin60;
        9'b000111101 : logsin3 = mux_in_sin61;
        9'b000111110 : logsin3 = mux_in_sin62;
        9'b000111111 : logsin3 = mux_in_sin63;
        9'b001000000 : logsin3 = mux_in_sin64;
        9'b001000001 : logsin3 = mux_in_sin65;
        9'b001000010 : logsin3 = mux_in_sin66;
        9'b001000011 : logsin3 = mux_in_sin67;
        9'b001000100 : logsin3 = mux_in_sin68;
        9'b001000101 : logsin3 = mux_in_sin69;
        9'b001000110 : logsin3 = mux_in_sin70;
        9'b001000111 : logsin3 = mux_in_sin71;
        9'b001001000 : logsin3 = mux_in_sin72;
        9'b001001001 : logsin3 = mux_in_sin73;
        9'b001001010 : logsin3 = mux_in_sin74;
        9'b001001011 : logsin3 = mux_in_sin75;
        9'b001001100 : logsin3 = mux_in_sin76;
        9'b001001101 : logsin3 = mux_in_sin77;
        9'b001001110 : logsin3 = mux_in_sin78;
        9'b001001111 : logsin3 = mux_in_sin79;
        9'b001010000 : logsin3 = mux_in_sin80;
        9'b001010001 : logsin3 = mux_in_sin81;
        9'b001010010 : logsin3 = mux_in_sin82;
        9'b001010011 : logsin3 = mux_in_sin83;
        9'b001010100 : logsin3 = mux_in_sin84;
        9'b001010101 : logsin3 = mux_in_sin85;
        9'b001010110 : logsin3 = mux_in_sin86;
        9'b001010111 : logsin3 = mux_in_sin87;
        9'b001011000 : logsin3 = mux_in_sin88;
        9'b001011001 : logsin3 = mux_in_sin89;
        9'b001011010 : logsin3 = mux_in_sin90;
        9'b001011011 : logsin3 = mux_in_sin91;
        9'b001011100 : logsin3 = mux_in_sin92;
        9'b001011101 : logsin3 = mux_in_sin93;
        9'b001011110 : logsin3 = mux_in_sin94;
        9'b001011111 : logsin3 = mux_in_sin95;
        9'b001100000 : logsin3 = mux_in_sin96;
        9'b001100001 : logsin3 = mux_in_sin97;
        9'b001100010 : logsin3 = mux_in_sin98;
        9'b001100011 : logsin3 = mux_in_sin99;
        9'b001100100 : logsin3 = mux_in_sin100;
        9'b001100101 : logsin3 = mux_in_sin101;
        9'b001100110 : logsin3 = mux_in_sin102;
        9'b001100111 : logsin3 = mux_in_sin103;
        9'b001101000 : logsin3 = mux_in_sin104;
        9'b001101001 : logsin3 = mux_in_sin105;
        9'b001101010 : logsin3 = mux_in_sin106;
        9'b001101011 : logsin3 = mux_in_sin107;
        9'b001101100 : logsin3 = mux_in_sin108;
        9'b001101101 : logsin3 = mux_in_sin109;
        9'b001101110 : logsin3 = mux_in_sin110;
        9'b001101111 : logsin3 = mux_in_sin111;
        9'b001110000 : logsin3 = mux_in_sin112;
        9'b001110001 : logsin3 = mux_in_sin113;
        9'b001110010 : logsin3 = mux_in_sin114;
        9'b001110011 : logsin3 = mux_in_sin115;
        9'b001110100 : logsin3 = mux_in_sin116;
        9'b001110101 : logsin3 = mux_in_sin117;
        9'b001110110 : logsin3 = mux_in_sin118;
        9'b001110111 : logsin3 = mux_in_sin119;
        9'b001111000 : logsin3 = mux_in_sin120;
        9'b001111001 : logsin3 = mux_in_sin121;
        9'b001111010 : logsin3 = mux_in_sin122;
        9'b001111011 : logsin3 = mux_in_sin123;
        9'b001111100 : logsin3 = mux_in_sin124;
        9'b001111101 : logsin3 = mux_in_sin125;
        9'b001111110 : logsin3 = mux_in_sin126;
        9'b001111111 : logsin3 = mux_in_sin127;
        9'b010000000 : logsin3 = mux_in_sin128;
        9'b010000001 : logsin3 = mux_in_sin129;
        9'b010000010 : logsin3 = mux_in_sin130;
        9'b010000011 : logsin3 = mux_in_sin131;
        9'b010000100 : logsin3 = mux_in_sin132;
        9'b010000101 : logsin3 = mux_in_sin133;
        9'b010000110 : logsin3 = mux_in_sin134;
        9'b010000111 : logsin3 = mux_in_sin135;
        9'b010001000 : logsin3 = mux_in_sin136;
        9'b010001001 : logsin3 = mux_in_sin137;
        9'b010001010 : logsin3 = mux_in_sin138;
        9'b010001011 : logsin3 = mux_in_sin139;
        9'b010001100 : logsin3 = mux_in_sin140;
        9'b010001101 : logsin3 = mux_in_sin141;
        9'b010001110 : logsin3 = mux_in_sin142;
        9'b010001111 : logsin3 = mux_in_sin143;
        9'b010010000 : logsin3 = mux_in_sin144;
        9'b010010001 : logsin3 = mux_in_sin145;
        9'b010010010 : logsin3 = mux_in_sin146;
        9'b010010011 : logsin3 = mux_in_sin147;
        9'b010010100 : logsin3 = mux_in_sin148;
        9'b010010101 : logsin3 = mux_in_sin149;
        9'b010010110 : logsin3 = mux_in_sin150;
        9'b010010111 : logsin3 = mux_in_sin151;
        9'b010011000 : logsin3 = mux_in_sin152;
        9'b010011001 : logsin3 = mux_in_sin153;
        9'b010011010 : logsin3 = mux_in_sin154;
        9'b010011011 : logsin3 = mux_in_sin155;
        9'b010011100 : logsin3 = mux_in_sin156;
        9'b010011101 : logsin3 = mux_in_sin157;
        9'b010011110 : logsin3 = mux_in_sin158;
        9'b010011111 : logsin3 = mux_in_sin159;
        9'b010100000 : logsin3 = mux_in_sin160;
        9'b010100001 : logsin3 = mux_in_sin161;
        9'b010100010 : logsin3 = mux_in_sin162;
        9'b010100011 : logsin3 = mux_in_sin163;
        9'b010100100 : logsin3 = mux_in_sin164;
        9'b010100101 : logsin3 = mux_in_sin165;
        9'b010100110 : logsin3 = mux_in_sin166;
        9'b010100111 : logsin3 = mux_in_sin167;
        9'b010101000 : logsin3 = mux_in_sin168;
        9'b010101001 : logsin3 = mux_in_sin169;
        9'b010101010 : logsin3 = mux_in_sin170;
        9'b010101011 : logsin3 = mux_in_sin171;
        9'b010101100 : logsin3 = mux_in_sin172;
        9'b010101101 : logsin3 = mux_in_sin173;
        9'b010101110 : logsin3 = mux_in_sin174;
        9'b010101111 : logsin3 = mux_in_sin175;
        9'b010110000 : logsin3 = mux_in_sin176;
        9'b010110001 : logsin3 = mux_in_sin177;
        9'b010110010 : logsin3 = mux_in_sin178;
        9'b010110011 : logsin3 = mux_in_sin179;
        9'b010110100 : logsin3 = mux_in_sin180;
        9'b010110101 : logsin3 = mux_in_sin181;
        9'b010110110 : logsin3 = mux_in_sin182;
        9'b010110111 : logsin3 = mux_in_sin183;
        9'b010111000 : logsin3 = mux_in_sin184;
        9'b010111001 : logsin3 = mux_in_sin185;
        9'b010111010 : logsin3 = mux_in_sin186;
        9'b010111011 : logsin3 = mux_in_sin187;
        9'b010111100 : logsin3 = mux_in_sin188;
        9'b010111101 : logsin3 = mux_in_sin189;
        9'b010111110 : logsin3 = mux_in_sin190;
        9'b010111111 : logsin3 = mux_in_sin191;
        9'b011000000 : logsin3 = mux_in_sin192;
        9'b011000001 : logsin3 = mux_in_sin193;
        9'b011000010 : logsin3 = mux_in_sin194;
        9'b011000011 : logsin3 = mux_in_sin195;
        9'b011000100 : logsin3 = mux_in_sin196;
        9'b011000101 : logsin3 = mux_in_sin197;
        9'b011000110 : logsin3 = mux_in_sin198;
        9'b011000111 : logsin3 = mux_in_sin199;
        9'b011001000 : logsin3 = mux_in_sin200;
        9'b011001001 : logsin3 = mux_in_sin201;
        9'b011001010 : logsin3 = mux_in_sin202;
        9'b011001011 : logsin3 = mux_in_sin203;
        9'b011001100 : logsin3 = mux_in_sin204;
        9'b011001101 : logsin3 = mux_in_sin205;
        9'b011001110 : logsin3 = mux_in_sin206;
        9'b011001111 : logsin3 = mux_in_sin207;
        9'b011010000 : logsin3 = mux_in_sin208;
        9'b011010001 : logsin3 = mux_in_sin209;
        9'b011010010 : logsin3 = mux_in_sin210;
        9'b011010011 : logsin3 = mux_in_sin211;
        9'b011010100 : logsin3 = mux_in_sin212;
        9'b011010101 : logsin3 = mux_in_sin213;
        9'b011010110 : logsin3 = mux_in_sin214;
        9'b011010111 : logsin3 = mux_in_sin215;
        9'b011011000 : logsin3 = mux_in_sin216;
        9'b011011001 : logsin3 = mux_in_sin217;
        9'b011011010 : logsin3 = mux_in_sin218;
        9'b011011011 : logsin3 = mux_in_sin219;
        9'b011011100 : logsin3 = mux_in_sin220;
        9'b011011101 : logsin3 = mux_in_sin221;
        9'b011011110 : logsin3 = mux_in_sin222;
        9'b011011111 : logsin3 = mux_in_sin223;
        9'b011100000 : logsin3 = mux_in_sin224;
        9'b011100001 : logsin3 = mux_in_sin225;
        9'b011100010 : logsin3 = mux_in_sin226;
        9'b011100011 : logsin3 = mux_in_sin227;
        9'b011100100 : logsin3 = mux_in_sin228;
        9'b011100101 : logsin3 = mux_in_sin229;
        9'b011100110 : logsin3 = mux_in_sin230;
        9'b011100111 : logsin3 = mux_in_sin231;
        9'b011101000 : logsin3 = mux_in_sin232;
        9'b011101001 : logsin3 = mux_in_sin233;
        9'b011101010 : logsin3 = mux_in_sin234;
        9'b011101011 : logsin3 = mux_in_sin235;
        9'b011101100 : logsin3 = mux_in_sin236;
        9'b011101101 : logsin3 = mux_in_sin237;
        9'b011101110 : logsin3 = mux_in_sin238;
        9'b011101111 : logsin3 = mux_in_sin239;
        9'b011110000 : logsin3 = mux_in_sin240;
        9'b011110001 : logsin3 = mux_in_sin241;
        9'b011110010 : logsin3 = mux_in_sin242;
        9'b011110011 : logsin3 = mux_in_sin243;
        9'b011110100 : logsin3 = mux_in_sin244;
        9'b011110101 : logsin3 = mux_in_sin245;
        9'b011110110 : logsin3 = mux_in_sin246;
        9'b011110111 : logsin3 = mux_in_sin247;
        9'b011111000 : logsin3 = mux_in_sin248;
        9'b011111001 : logsin3 = mux_in_sin249;
        9'b011111010 : logsin3 = mux_in_sin250;
        9'b011111011 : logsin3 = mux_in_sin251;
        9'b011111100 : logsin3 = mux_in_sin252;
        9'b011111101 : logsin3 = mux_in_sin253;
        9'b011111110 : logsin3 = mux_in_sin254;
        9'b011111111 : logsin3 = mux_in_sin255;
        9'b100000000 : logsin3 = mux_in_sin256;
        default: logsin3 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in1)
        9'b000000000 : logcos1 = mux_in_cos0;
        9'b000000001 : logcos1 = mux_in_cos1;
        9'b000000010 : logcos1 = mux_in_cos2;
        9'b000000011 : logcos1 = mux_in_cos3;
        9'b000000100 : logcos1 = mux_in_cos4;
        9'b000000101 : logcos1 = mux_in_cos5;
        9'b000000110 : logcos1 = mux_in_cos6;
        9'b000000111 : logcos1 = mux_in_cos7;
        9'b000001000 : logcos1 = mux_in_cos8;
        9'b000001001 : logcos1 = mux_in_cos9;
        9'b000001010 : logcos1 = mux_in_cos10;
        9'b000001011 : logcos1 = mux_in_cos11;
        9'b000001100 : logcos1 = mux_in_cos12;
        9'b000001101 : logcos1 = mux_in_cos13;
        9'b000001110 : logcos1 = mux_in_cos14;
        9'b000001111 : logcos1 = mux_in_cos15;
        9'b000010000 : logcos1 = mux_in_cos16;
        9'b000010001 : logcos1 = mux_in_cos17;
        9'b000010010 : logcos1 = mux_in_cos18;
        9'b000010011 : logcos1 = mux_in_cos19;
        9'b000010100 : logcos1 = mux_in_cos20;
        9'b000010101 : logcos1 = mux_in_cos21;
        9'b000010110 : logcos1 = mux_in_cos22;
        9'b000010111 : logcos1 = mux_in_cos23;
        9'b000011000 : logcos1 = mux_in_cos24;
        9'b000011001 : logcos1 = mux_in_cos25;
        9'b000011010 : logcos1 = mux_in_cos26;
        9'b000011011 : logcos1 = mux_in_cos27;
        9'b000011100 : logcos1 = mux_in_cos28;
        9'b000011101 : logcos1 = mux_in_cos29;
        9'b000011110 : logcos1 = mux_in_cos30;
        9'b000011111 : logcos1 = mux_in_cos31;
        9'b000100000 : logcos1 = mux_in_cos32;
        9'b000100001 : logcos1 = mux_in_cos33;
        9'b000100010 : logcos1 = mux_in_cos34;
        9'b000100011 : logcos1 = mux_in_cos35;
        9'b000100100 : logcos1 = mux_in_cos36;
        9'b000100101 : logcos1 = mux_in_cos37;
        9'b000100110 : logcos1 = mux_in_cos38;
        9'b000100111 : logcos1 = mux_in_cos39;
        9'b000101000 : logcos1 = mux_in_cos40;
        9'b000101001 : logcos1 = mux_in_cos41;
        9'b000101010 : logcos1 = mux_in_cos42;
        9'b000101011 : logcos1 = mux_in_cos43;
        9'b000101100 : logcos1 = mux_in_cos44;
        9'b000101101 : logcos1 = mux_in_cos45;
        9'b000101110 : logcos1 = mux_in_cos46;
        9'b000101111 : logcos1 = mux_in_cos47;
        9'b000110000 : logcos1 = mux_in_cos48;
        9'b000110001 : logcos1 = mux_in_cos49;
        9'b000110010 : logcos1 = mux_in_cos50;
        9'b000110011 : logcos1 = mux_in_cos51;
        9'b000110100 : logcos1 = mux_in_cos52;
        9'b000110101 : logcos1 = mux_in_cos53;
        9'b000110110 : logcos1 = mux_in_cos54;
        9'b000110111 : logcos1 = mux_in_cos55;
        9'b000111000 : logcos1 = mux_in_cos56;
        9'b000111001 : logcos1 = mux_in_cos57;
        9'b000111010 : logcos1 = mux_in_cos58;
        9'b000111011 : logcos1 = mux_in_cos59;
        9'b000111100 : logcos1 = mux_in_cos60;
        9'b000111101 : logcos1 = mux_in_cos61;
        9'b000111110 : logcos1 = mux_in_cos62;
        9'b000111111 : logcos1 = mux_in_cos63;
        9'b001000000 : logcos1 = mux_in_cos64;
        9'b001000001 : logcos1 = mux_in_cos65;
        9'b001000010 : logcos1 = mux_in_cos66;
        9'b001000011 : logcos1 = mux_in_cos67;
        9'b001000100 : logcos1 = mux_in_cos68;
        9'b001000101 : logcos1 = mux_in_cos69;
        9'b001000110 : logcos1 = mux_in_cos70;
        9'b001000111 : logcos1 = mux_in_cos71;
        9'b001001000 : logcos1 = mux_in_cos72;
        9'b001001001 : logcos1 = mux_in_cos73;
        9'b001001010 : logcos1 = mux_in_cos74;
        9'b001001011 : logcos1 = mux_in_cos75;
        9'b001001100 : logcos1 = mux_in_cos76;
        9'b001001101 : logcos1 = mux_in_cos77;
        9'b001001110 : logcos1 = mux_in_cos78;
        9'b001001111 : logcos1 = mux_in_cos79;
        9'b001010000 : logcos1 = mux_in_cos80;
        9'b001010001 : logcos1 = mux_in_cos81;
        9'b001010010 : logcos1 = mux_in_cos82;
        9'b001010011 : logcos1 = mux_in_cos83;
        9'b001010100 : logcos1 = mux_in_cos84;
        9'b001010101 : logcos1 = mux_in_cos85;
        9'b001010110 : logcos1 = mux_in_cos86;
        9'b001010111 : logcos1 = mux_in_cos87;
        9'b001011000 : logcos1 = mux_in_cos88;
        9'b001011001 : logcos1 = mux_in_cos89;
        9'b001011010 : logcos1 = mux_in_cos90;
        9'b001011011 : logcos1 = mux_in_cos91;
        9'b001011100 : logcos1 = mux_in_cos92;
        9'b001011101 : logcos1 = mux_in_cos93;
        9'b001011110 : logcos1 = mux_in_cos94;
        9'b001011111 : logcos1 = mux_in_cos95;
        9'b001100000 : logcos1 = mux_in_cos96;
        9'b001100001 : logcos1 = mux_in_cos97;
        9'b001100010 : logcos1 = mux_in_cos98;
        9'b001100011 : logcos1 = mux_in_cos99;
        9'b001100100 : logcos1 = mux_in_cos100;
        9'b001100101 : logcos1 = mux_in_cos101;
        9'b001100110 : logcos1 = mux_in_cos102;
        9'b001100111 : logcos1 = mux_in_cos103;
        9'b001101000 : logcos1 = mux_in_cos104;
        9'b001101001 : logcos1 = mux_in_cos105;
        9'b001101010 : logcos1 = mux_in_cos106;
        9'b001101011 : logcos1 = mux_in_cos107;
        9'b001101100 : logcos1 = mux_in_cos108;
        9'b001101101 : logcos1 = mux_in_cos109;
        9'b001101110 : logcos1 = mux_in_cos110;
        9'b001101111 : logcos1 = mux_in_cos111;
        9'b001110000 : logcos1 = mux_in_cos112;
        9'b001110001 : logcos1 = mux_in_cos113;
        9'b001110010 : logcos1 = mux_in_cos114;
        9'b001110011 : logcos1 = mux_in_cos115;
        9'b001110100 : logcos1 = mux_in_cos116;
        9'b001110101 : logcos1 = mux_in_cos117;
        9'b001110110 : logcos1 = mux_in_cos118;
        9'b001110111 : logcos1 = mux_in_cos119;
        9'b001111000 : logcos1 = mux_in_cos120;
        9'b001111001 : logcos1 = mux_in_cos121;
        9'b001111010 : logcos1 = mux_in_cos122;
        9'b001111011 : logcos1 = mux_in_cos123;
        9'b001111100 : logcos1 = mux_in_cos124;
        9'b001111101 : logcos1 = mux_in_cos125;
        9'b001111110 : logcos1 = mux_in_cos126;
        9'b001111111 : logcos1 = mux_in_cos127;
        9'b010000000 : logcos1 = mux_in_cos128;
        9'b010000001 : logcos1 = mux_in_cos129;
        9'b010000010 : logcos1 = mux_in_cos130;
        9'b010000011 : logcos1 = mux_in_cos131;
        9'b010000100 : logcos1 = mux_in_cos132;
        9'b010000101 : logcos1 = mux_in_cos133;
        9'b010000110 : logcos1 = mux_in_cos134;
        9'b010000111 : logcos1 = mux_in_cos135;
        9'b010001000 : logcos1 = mux_in_cos136;
        9'b010001001 : logcos1 = mux_in_cos137;
        9'b010001010 : logcos1 = mux_in_cos138;
        9'b010001011 : logcos1 = mux_in_cos139;
        9'b010001100 : logcos1 = mux_in_cos140;
        9'b010001101 : logcos1 = mux_in_cos141;
        9'b010001110 : logcos1 = mux_in_cos142;
        9'b010001111 : logcos1 = mux_in_cos143;
        9'b010010000 : logcos1 = mux_in_cos144;
        9'b010010001 : logcos1 = mux_in_cos145;
        9'b010010010 : logcos1 = mux_in_cos146;
        9'b010010011 : logcos1 = mux_in_cos147;
        9'b010010100 : logcos1 = mux_in_cos148;
        9'b010010101 : logcos1 = mux_in_cos149;
        9'b010010110 : logcos1 = mux_in_cos150;
        9'b010010111 : logcos1 = mux_in_cos151;
        9'b010011000 : logcos1 = mux_in_cos152;
        9'b010011001 : logcos1 = mux_in_cos153;
        9'b010011010 : logcos1 = mux_in_cos154;
        9'b010011011 : logcos1 = mux_in_cos155;
        9'b010011100 : logcos1 = mux_in_cos156;
        9'b010011101 : logcos1 = mux_in_cos157;
        9'b010011110 : logcos1 = mux_in_cos158;
        9'b010011111 : logcos1 = mux_in_cos159;
        9'b010100000 : logcos1 = mux_in_cos160;
        9'b010100001 : logcos1 = mux_in_cos161;
        9'b010100010 : logcos1 = mux_in_cos162;
        9'b010100011 : logcos1 = mux_in_cos163;
        9'b010100100 : logcos1 = mux_in_cos164;
        9'b010100101 : logcos1 = mux_in_cos165;
        9'b010100110 : logcos1 = mux_in_cos166;
        9'b010100111 : logcos1 = mux_in_cos167;
        9'b010101000 : logcos1 = mux_in_cos168;
        9'b010101001 : logcos1 = mux_in_cos169;
        9'b010101010 : logcos1 = mux_in_cos170;
        9'b010101011 : logcos1 = mux_in_cos171;
        9'b010101100 : logcos1 = mux_in_cos172;
        9'b010101101 : logcos1 = mux_in_cos173;
        9'b010101110 : logcos1 = mux_in_cos174;
        9'b010101111 : logcos1 = mux_in_cos175;
        9'b010110000 : logcos1 = mux_in_cos176;
        9'b010110001 : logcos1 = mux_in_cos177;
        9'b010110010 : logcos1 = mux_in_cos178;
        9'b010110011 : logcos1 = mux_in_cos179;
        9'b010110100 : logcos1 = mux_in_cos180;
        9'b010110101 : logcos1 = mux_in_cos181;
        9'b010110110 : logcos1 = mux_in_cos182;
        9'b010110111 : logcos1 = mux_in_cos183;
        9'b010111000 : logcos1 = mux_in_cos184;
        9'b010111001 : logcos1 = mux_in_cos185;
        9'b010111010 : logcos1 = mux_in_cos186;
        9'b010111011 : logcos1 = mux_in_cos187;
        9'b010111100 : logcos1 = mux_in_cos188;
        9'b010111101 : logcos1 = mux_in_cos189;
        9'b010111110 : logcos1 = mux_in_cos190;
        9'b010111111 : logcos1 = mux_in_cos191;
        9'b011000000 : logcos1 = mux_in_cos192;
        9'b011000001 : logcos1 = mux_in_cos193;
        9'b011000010 : logcos1 = mux_in_cos194;
        9'b011000011 : logcos1 = mux_in_cos195;
        9'b011000100 : logcos1 = mux_in_cos196;
        9'b011000101 : logcos1 = mux_in_cos197;
        9'b011000110 : logcos1 = mux_in_cos198;
        9'b011000111 : logcos1 = mux_in_cos199;
        9'b011001000 : logcos1 = mux_in_cos200;
        9'b011001001 : logcos1 = mux_in_cos201;
        9'b011001010 : logcos1 = mux_in_cos202;
        9'b011001011 : logcos1 = mux_in_cos203;
        9'b011001100 : logcos1 = mux_in_cos204;
        9'b011001101 : logcos1 = mux_in_cos205;
        9'b011001110 : logcos1 = mux_in_cos206;
        9'b011001111 : logcos1 = mux_in_cos207;
        9'b011010000 : logcos1 = mux_in_cos208;
        9'b011010001 : logcos1 = mux_in_cos209;
        9'b011010010 : logcos1 = mux_in_cos210;
        9'b011010011 : logcos1 = mux_in_cos211;
        9'b011010100 : logcos1 = mux_in_cos212;
        9'b011010101 : logcos1 = mux_in_cos213;
        9'b011010110 : logcos1 = mux_in_cos214;
        9'b011010111 : logcos1 = mux_in_cos215;
        9'b011011000 : logcos1 = mux_in_cos216;
        9'b011011001 : logcos1 = mux_in_cos217;
        9'b011011010 : logcos1 = mux_in_cos218;
        9'b011011011 : logcos1 = mux_in_cos219;
        9'b011011100 : logcos1 = mux_in_cos220;
        9'b011011101 : logcos1 = mux_in_cos221;
        9'b011011110 : logcos1 = mux_in_cos222;
        9'b011011111 : logcos1 = mux_in_cos223;
        9'b011100000 : logcos1 = mux_in_cos224;
        9'b011100001 : logcos1 = mux_in_cos225;
        9'b011100010 : logcos1 = mux_in_cos226;
        9'b011100011 : logcos1 = mux_in_cos227;
        9'b011100100 : logcos1 = mux_in_cos228;
        9'b011100101 : logcos1 = mux_in_cos229;
        9'b011100110 : logcos1 = mux_in_cos230;
        9'b011100111 : logcos1 = mux_in_cos231;
        9'b011101000 : logcos1 = mux_in_cos232;
        9'b011101001 : logcos1 = mux_in_cos233;
        9'b011101010 : logcos1 = mux_in_cos234;
        9'b011101011 : logcos1 = mux_in_cos235;
        9'b011101100 : logcos1 = mux_in_cos236;
        9'b011101101 : logcos1 = mux_in_cos237;
        9'b011101110 : logcos1 = mux_in_cos238;
        9'b011101111 : logcos1 = mux_in_cos239;
        9'b011110000 : logcos1 = mux_in_cos240;
        9'b011110001 : logcos1 = mux_in_cos241;
        9'b011110010 : logcos1 = mux_in_cos242;
        9'b011110011 : logcos1 = mux_in_cos243;
        9'b011110100 : logcos1 = mux_in_cos244;
        9'b011110101 : logcos1 = mux_in_cos245;
        9'b011110110 : logcos1 = mux_in_cos246;
        9'b011110111 : logcos1 = mux_in_cos247;
        9'b011111000 : logcos1 = mux_in_cos248;
        9'b011111001 : logcos1 = mux_in_cos249;
        9'b011111010 : logcos1 = mux_in_cos250;
        9'b011111011 : logcos1 = mux_in_cos251;
        9'b011111100 : logcos1 = mux_in_cos252;
        9'b011111101 : logcos1 = mux_in_cos253;
        9'b011111110 : logcos1 = mux_in_cos254;
        9'b011111111 : logcos1 = mux_in_cos255;
        9'b100000000 : logcos1 = mux_in_cos256;
        default: logcos1 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in2)
        9'b000000000 : logcos2 = mux_in_cos0;
        9'b000000001 : logcos2 = mux_in_cos1;
        9'b000000010 : logcos2 = mux_in_cos2;
        9'b000000011 : logcos2 = mux_in_cos3;
        9'b000000100 : logcos2 = mux_in_cos4;
        9'b000000101 : logcos2 = mux_in_cos5;
        9'b000000110 : logcos2 = mux_in_cos6;
        9'b000000111 : logcos2 = mux_in_cos7;
        9'b000001000 : logcos2 = mux_in_cos8;
        9'b000001001 : logcos2 = mux_in_cos9;
        9'b000001010 : logcos2 = mux_in_cos10;
        9'b000001011 : logcos2 = mux_in_cos11;
        9'b000001100 : logcos2 = mux_in_cos12;
        9'b000001101 : logcos2 = mux_in_cos13;
        9'b000001110 : logcos2 = mux_in_cos14;
        9'b000001111 : logcos2 = mux_in_cos15;
        9'b000010000 : logcos2 = mux_in_cos16;
        9'b000010001 : logcos2 = mux_in_cos17;
        9'b000010010 : logcos2 = mux_in_cos18;
        9'b000010011 : logcos2 = mux_in_cos19;
        9'b000010100 : logcos2 = mux_in_cos20;
        9'b000010101 : logcos2 = mux_in_cos21;
        9'b000010110 : logcos2 = mux_in_cos22;
        9'b000010111 : logcos2 = mux_in_cos23;
        9'b000011000 : logcos2 = mux_in_cos24;
        9'b000011001 : logcos2 = mux_in_cos25;
        9'b000011010 : logcos2 = mux_in_cos26;
        9'b000011011 : logcos2 = mux_in_cos27;
        9'b000011100 : logcos2 = mux_in_cos28;
        9'b000011101 : logcos2 = mux_in_cos29;
        9'b000011110 : logcos2 = mux_in_cos30;
        9'b000011111 : logcos2 = mux_in_cos31;
        9'b000100000 : logcos2 = mux_in_cos32;
        9'b000100001 : logcos2 = mux_in_cos33;
        9'b000100010 : logcos2 = mux_in_cos34;
        9'b000100011 : logcos2 = mux_in_cos35;
        9'b000100100 : logcos2 = mux_in_cos36;
        9'b000100101 : logcos2 = mux_in_cos37;
        9'b000100110 : logcos2 = mux_in_cos38;
        9'b000100111 : logcos2 = mux_in_cos39;
        9'b000101000 : logcos2 = mux_in_cos40;
        9'b000101001 : logcos2 = mux_in_cos41;
        9'b000101010 : logcos2 = mux_in_cos42;
        9'b000101011 : logcos2 = mux_in_cos43;
        9'b000101100 : logcos2 = mux_in_cos44;
        9'b000101101 : logcos2 = mux_in_cos45;
        9'b000101110 : logcos2 = mux_in_cos46;
        9'b000101111 : logcos2 = mux_in_cos47;
        9'b000110000 : logcos2 = mux_in_cos48;
        9'b000110001 : logcos2 = mux_in_cos49;
        9'b000110010 : logcos2 = mux_in_cos50;
        9'b000110011 : logcos2 = mux_in_cos51;
        9'b000110100 : logcos2 = mux_in_cos52;
        9'b000110101 : logcos2 = mux_in_cos53;
        9'b000110110 : logcos2 = mux_in_cos54;
        9'b000110111 : logcos2 = mux_in_cos55;
        9'b000111000 : logcos2 = mux_in_cos56;
        9'b000111001 : logcos2 = mux_in_cos57;
        9'b000111010 : logcos2 = mux_in_cos58;
        9'b000111011 : logcos2 = mux_in_cos59;
        9'b000111100 : logcos2 = mux_in_cos60;
        9'b000111101 : logcos2 = mux_in_cos61;
        9'b000111110 : logcos2 = mux_in_cos62;
        9'b000111111 : logcos2 = mux_in_cos63;
        9'b001000000 : logcos2 = mux_in_cos64;
        9'b001000001 : logcos2 = mux_in_cos65;
        9'b001000010 : logcos2 = mux_in_cos66;
        9'b001000011 : logcos2 = mux_in_cos67;
        9'b001000100 : logcos2 = mux_in_cos68;
        9'b001000101 : logcos2 = mux_in_cos69;
        9'b001000110 : logcos2 = mux_in_cos70;
        9'b001000111 : logcos2 = mux_in_cos71;
        9'b001001000 : logcos2 = mux_in_cos72;
        9'b001001001 : logcos2 = mux_in_cos73;
        9'b001001010 : logcos2 = mux_in_cos74;
        9'b001001011 : logcos2 = mux_in_cos75;
        9'b001001100 : logcos2 = mux_in_cos76;
        9'b001001101 : logcos2 = mux_in_cos77;
        9'b001001110 : logcos2 = mux_in_cos78;
        9'b001001111 : logcos2 = mux_in_cos79;
        9'b001010000 : logcos2 = mux_in_cos80;
        9'b001010001 : logcos2 = mux_in_cos81;
        9'b001010010 : logcos2 = mux_in_cos82;
        9'b001010011 : logcos2 = mux_in_cos83;
        9'b001010100 : logcos2 = mux_in_cos84;
        9'b001010101 : logcos2 = mux_in_cos85;
        9'b001010110 : logcos2 = mux_in_cos86;
        9'b001010111 : logcos2 = mux_in_cos87;
        9'b001011000 : logcos2 = mux_in_cos88;
        9'b001011001 : logcos2 = mux_in_cos89;
        9'b001011010 : logcos2 = mux_in_cos90;
        9'b001011011 : logcos2 = mux_in_cos91;
        9'b001011100 : logcos2 = mux_in_cos92;
        9'b001011101 : logcos2 = mux_in_cos93;
        9'b001011110 : logcos2 = mux_in_cos94;
        9'b001011111 : logcos2 = mux_in_cos95;
        9'b001100000 : logcos2 = mux_in_cos96;
        9'b001100001 : logcos2 = mux_in_cos97;
        9'b001100010 : logcos2 = mux_in_cos98;
        9'b001100011 : logcos2 = mux_in_cos99;
        9'b001100100 : logcos2 = mux_in_cos100;
        9'b001100101 : logcos2 = mux_in_cos101;
        9'b001100110 : logcos2 = mux_in_cos102;
        9'b001100111 : logcos2 = mux_in_cos103;
        9'b001101000 : logcos2 = mux_in_cos104;
        9'b001101001 : logcos2 = mux_in_cos105;
        9'b001101010 : logcos2 = mux_in_cos106;
        9'b001101011 : logcos2 = mux_in_cos107;
        9'b001101100 : logcos2 = mux_in_cos108;
        9'b001101101 : logcos2 = mux_in_cos109;
        9'b001101110 : logcos2 = mux_in_cos110;
        9'b001101111 : logcos2 = mux_in_cos111;
        9'b001110000 : logcos2 = mux_in_cos112;
        9'b001110001 : logcos2 = mux_in_cos113;
        9'b001110010 : logcos2 = mux_in_cos114;
        9'b001110011 : logcos2 = mux_in_cos115;
        9'b001110100 : logcos2 = mux_in_cos116;
        9'b001110101 : logcos2 = mux_in_cos117;
        9'b001110110 : logcos2 = mux_in_cos118;
        9'b001110111 : logcos2 = mux_in_cos119;
        9'b001111000 : logcos2 = mux_in_cos120;
        9'b001111001 : logcos2 = mux_in_cos121;
        9'b001111010 : logcos2 = mux_in_cos122;
        9'b001111011 : logcos2 = mux_in_cos123;
        9'b001111100 : logcos2 = mux_in_cos124;
        9'b001111101 : logcos2 = mux_in_cos125;
        9'b001111110 : logcos2 = mux_in_cos126;
        9'b001111111 : logcos2 = mux_in_cos127;
        9'b010000000 : logcos2 = mux_in_cos128;
        9'b010000001 : logcos2 = mux_in_cos129;
        9'b010000010 : logcos2 = mux_in_cos130;
        9'b010000011 : logcos2 = mux_in_cos131;
        9'b010000100 : logcos2 = mux_in_cos132;
        9'b010000101 : logcos2 = mux_in_cos133;
        9'b010000110 : logcos2 = mux_in_cos134;
        9'b010000111 : logcos2 = mux_in_cos135;
        9'b010001000 : logcos2 = mux_in_cos136;
        9'b010001001 : logcos2 = mux_in_cos137;
        9'b010001010 : logcos2 = mux_in_cos138;
        9'b010001011 : logcos2 = mux_in_cos139;
        9'b010001100 : logcos2 = mux_in_cos140;
        9'b010001101 : logcos2 = mux_in_cos141;
        9'b010001110 : logcos2 = mux_in_cos142;
        9'b010001111 : logcos2 = mux_in_cos143;
        9'b010010000 : logcos2 = mux_in_cos144;
        9'b010010001 : logcos2 = mux_in_cos145;
        9'b010010010 : logcos2 = mux_in_cos146;
        9'b010010011 : logcos2 = mux_in_cos147;
        9'b010010100 : logcos2 = mux_in_cos148;
        9'b010010101 : logcos2 = mux_in_cos149;
        9'b010010110 : logcos2 = mux_in_cos150;
        9'b010010111 : logcos2 = mux_in_cos151;
        9'b010011000 : logcos2 = mux_in_cos152;
        9'b010011001 : logcos2 = mux_in_cos153;
        9'b010011010 : logcos2 = mux_in_cos154;
        9'b010011011 : logcos2 = mux_in_cos155;
        9'b010011100 : logcos2 = mux_in_cos156;
        9'b010011101 : logcos2 = mux_in_cos157;
        9'b010011110 : logcos2 = mux_in_cos158;
        9'b010011111 : logcos2 = mux_in_cos159;
        9'b010100000 : logcos2 = mux_in_cos160;
        9'b010100001 : logcos2 = mux_in_cos161;
        9'b010100010 : logcos2 = mux_in_cos162;
        9'b010100011 : logcos2 = mux_in_cos163;
        9'b010100100 : logcos2 = mux_in_cos164;
        9'b010100101 : logcos2 = mux_in_cos165;
        9'b010100110 : logcos2 = mux_in_cos166;
        9'b010100111 : logcos2 = mux_in_cos167;
        9'b010101000 : logcos2 = mux_in_cos168;
        9'b010101001 : logcos2 = mux_in_cos169;
        9'b010101010 : logcos2 = mux_in_cos170;
        9'b010101011 : logcos2 = mux_in_cos171;
        9'b010101100 : logcos2 = mux_in_cos172;
        9'b010101101 : logcos2 = mux_in_cos173;
        9'b010101110 : logcos2 = mux_in_cos174;
        9'b010101111 : logcos2 = mux_in_cos175;
        9'b010110000 : logcos2 = mux_in_cos176;
        9'b010110001 : logcos2 = mux_in_cos177;
        9'b010110010 : logcos2 = mux_in_cos178;
        9'b010110011 : logcos2 = mux_in_cos179;
        9'b010110100 : logcos2 = mux_in_cos180;
        9'b010110101 : logcos2 = mux_in_cos181;
        9'b010110110 : logcos2 = mux_in_cos182;
        9'b010110111 : logcos2 = mux_in_cos183;
        9'b010111000 : logcos2 = mux_in_cos184;
        9'b010111001 : logcos2 = mux_in_cos185;
        9'b010111010 : logcos2 = mux_in_cos186;
        9'b010111011 : logcos2 = mux_in_cos187;
        9'b010111100 : logcos2 = mux_in_cos188;
        9'b010111101 : logcos2 = mux_in_cos189;
        9'b010111110 : logcos2 = mux_in_cos190;
        9'b010111111 : logcos2 = mux_in_cos191;
        9'b011000000 : logcos2 = mux_in_cos192;
        9'b011000001 : logcos2 = mux_in_cos193;
        9'b011000010 : logcos2 = mux_in_cos194;
        9'b011000011 : logcos2 = mux_in_cos195;
        9'b011000100 : logcos2 = mux_in_cos196;
        9'b011000101 : logcos2 = mux_in_cos197;
        9'b011000110 : logcos2 = mux_in_cos198;
        9'b011000111 : logcos2 = mux_in_cos199;
        9'b011001000 : logcos2 = mux_in_cos200;
        9'b011001001 : logcos2 = mux_in_cos201;
        9'b011001010 : logcos2 = mux_in_cos202;
        9'b011001011 : logcos2 = mux_in_cos203;
        9'b011001100 : logcos2 = mux_in_cos204;
        9'b011001101 : logcos2 = mux_in_cos205;
        9'b011001110 : logcos2 = mux_in_cos206;
        9'b011001111 : logcos2 = mux_in_cos207;
        9'b011010000 : logcos2 = mux_in_cos208;
        9'b011010001 : logcos2 = mux_in_cos209;
        9'b011010010 : logcos2 = mux_in_cos210;
        9'b011010011 : logcos2 = mux_in_cos211;
        9'b011010100 : logcos2 = mux_in_cos212;
        9'b011010101 : logcos2 = mux_in_cos213;
        9'b011010110 : logcos2 = mux_in_cos214;
        9'b011010111 : logcos2 = mux_in_cos215;
        9'b011011000 : logcos2 = mux_in_cos216;
        9'b011011001 : logcos2 = mux_in_cos217;
        9'b011011010 : logcos2 = mux_in_cos218;
        9'b011011011 : logcos2 = mux_in_cos219;
        9'b011011100 : logcos2 = mux_in_cos220;
        9'b011011101 : logcos2 = mux_in_cos221;
        9'b011011110 : logcos2 = mux_in_cos222;
        9'b011011111 : logcos2 = mux_in_cos223;
        9'b011100000 : logcos2 = mux_in_cos224;
        9'b011100001 : logcos2 = mux_in_cos225;
        9'b011100010 : logcos2 = mux_in_cos226;
        9'b011100011 : logcos2 = mux_in_cos227;
        9'b011100100 : logcos2 = mux_in_cos228;
        9'b011100101 : logcos2 = mux_in_cos229;
        9'b011100110 : logcos2 = mux_in_cos230;
        9'b011100111 : logcos2 = mux_in_cos231;
        9'b011101000 : logcos2 = mux_in_cos232;
        9'b011101001 : logcos2 = mux_in_cos233;
        9'b011101010 : logcos2 = mux_in_cos234;
        9'b011101011 : logcos2 = mux_in_cos235;
        9'b011101100 : logcos2 = mux_in_cos236;
        9'b011101101 : logcos2 = mux_in_cos237;
        9'b011101110 : logcos2 = mux_in_cos238;
        9'b011101111 : logcos2 = mux_in_cos239;
        9'b011110000 : logcos2 = mux_in_cos240;
        9'b011110001 : logcos2 = mux_in_cos241;
        9'b011110010 : logcos2 = mux_in_cos242;
        9'b011110011 : logcos2 = mux_in_cos243;
        9'b011110100 : logcos2 = mux_in_cos244;
        9'b011110101 : logcos2 = mux_in_cos245;
        9'b011110110 : logcos2 = mux_in_cos246;
        9'b011110111 : logcos2 = mux_in_cos247;
        9'b011111000 : logcos2 = mux_in_cos248;
        9'b011111001 : logcos2 = mux_in_cos249;
        9'b011111010 : logcos2 = mux_in_cos250;
        9'b011111011 : logcos2 = mux_in_cos251;
        9'b011111100 : logcos2 = mux_in_cos252;
        9'b011111101 : logcos2 = mux_in_cos253;
        9'b011111110 : logcos2 = mux_in_cos254;
        9'b011111111 : logcos2 = mux_in_cos255;
        9'b100000000 : logcos2 = mux_in_cos256;
        default: logcos2 = 15'bx;
        endcase
    end

    always @ (*)
    begin
        case(x_in3)
        9'b000000000 : logcos3 = mux_in_cos0;
        9'b000000001 : logcos3 = mux_in_cos1;
        9'b000000010 : logcos3 = mux_in_cos2;
        9'b000000011 : logcos3 = mux_in_cos3;
        9'b000000100 : logcos3 = mux_in_cos4;
        9'b000000101 : logcos3 = mux_in_cos5;
        9'b000000110 : logcos3 = mux_in_cos6;
        9'b000000111 : logcos3 = mux_in_cos7;
        9'b000001000 : logcos3 = mux_in_cos8;
        9'b000001001 : logcos3 = mux_in_cos9;
        9'b000001010 : logcos3 = mux_in_cos10;
        9'b000001011 : logcos3 = mux_in_cos11;
        9'b000001100 : logcos3 = mux_in_cos12;
        9'b000001101 : logcos3 = mux_in_cos13;
        9'b000001110 : logcos3 = mux_in_cos14;
        9'b000001111 : logcos3 = mux_in_cos15;
        9'b000010000 : logcos3 = mux_in_cos16;
        9'b000010001 : logcos3 = mux_in_cos17;
        9'b000010010 : logcos3 = mux_in_cos18;
        9'b000010011 : logcos3 = mux_in_cos19;
        9'b000010100 : logcos3 = mux_in_cos20;
        9'b000010101 : logcos3 = mux_in_cos21;
        9'b000010110 : logcos3 = mux_in_cos22;
        9'b000010111 : logcos3 = mux_in_cos23;
        9'b000011000 : logcos3 = mux_in_cos24;
        9'b000011001 : logcos3 = mux_in_cos25;
        9'b000011010 : logcos3 = mux_in_cos26;
        9'b000011011 : logcos3 = mux_in_cos27;
        9'b000011100 : logcos3 = mux_in_cos28;
        9'b000011101 : logcos3 = mux_in_cos29;
        9'b000011110 : logcos3 = mux_in_cos30;
        9'b000011111 : logcos3 = mux_in_cos31;
        9'b000100000 : logcos3 = mux_in_cos32;
        9'b000100001 : logcos3 = mux_in_cos33;
        9'b000100010 : logcos3 = mux_in_cos34;
        9'b000100011 : logcos3 = mux_in_cos35;
        9'b000100100 : logcos3 = mux_in_cos36;
        9'b000100101 : logcos3 = mux_in_cos37;
        9'b000100110 : logcos3 = mux_in_cos38;
        9'b000100111 : logcos3 = mux_in_cos39;
        9'b000101000 : logcos3 = mux_in_cos40;
        9'b000101001 : logcos3 = mux_in_cos41;
        9'b000101010 : logcos3 = mux_in_cos42;
        9'b000101011 : logcos3 = mux_in_cos43;
        9'b000101100 : logcos3 = mux_in_cos44;
        9'b000101101 : logcos3 = mux_in_cos45;
        9'b000101110 : logcos3 = mux_in_cos46;
        9'b000101111 : logcos3 = mux_in_cos47;
        9'b000110000 : logcos3 = mux_in_cos48;
        9'b000110001 : logcos3 = mux_in_cos49;
        9'b000110010 : logcos3 = mux_in_cos50;
        9'b000110011 : logcos3 = mux_in_cos51;
        9'b000110100 : logcos3 = mux_in_cos52;
        9'b000110101 : logcos3 = mux_in_cos53;
        9'b000110110 : logcos3 = mux_in_cos54;
        9'b000110111 : logcos3 = mux_in_cos55;
        9'b000111000 : logcos3 = mux_in_cos56;
        9'b000111001 : logcos3 = mux_in_cos57;
        9'b000111010 : logcos3 = mux_in_cos58;
        9'b000111011 : logcos3 = mux_in_cos59;
        9'b000111100 : logcos3 = mux_in_cos60;
        9'b000111101 : logcos3 = mux_in_cos61;
        9'b000111110 : logcos3 = mux_in_cos62;
        9'b000111111 : logcos3 = mux_in_cos63;
        9'b001000000 : logcos3 = mux_in_cos64;
        9'b001000001 : logcos3 = mux_in_cos65;
        9'b001000010 : logcos3 = mux_in_cos66;
        9'b001000011 : logcos3 = mux_in_cos67;
        9'b001000100 : logcos3 = mux_in_cos68;
        9'b001000101 : logcos3 = mux_in_cos69;
        9'b001000110 : logcos3 = mux_in_cos70;
        9'b001000111 : logcos3 = mux_in_cos71;
        9'b001001000 : logcos3 = mux_in_cos72;
        9'b001001001 : logcos3 = mux_in_cos73;
        9'b001001010 : logcos3 = mux_in_cos74;
        9'b001001011 : logcos3 = mux_in_cos75;
        9'b001001100 : logcos3 = mux_in_cos76;
        9'b001001101 : logcos3 = mux_in_cos77;
        9'b001001110 : logcos3 = mux_in_cos78;
        9'b001001111 : logcos3 = mux_in_cos79;
        9'b001010000 : logcos3 = mux_in_cos80;
        9'b001010001 : logcos3 = mux_in_cos81;
        9'b001010010 : logcos3 = mux_in_cos82;
        9'b001010011 : logcos3 = mux_in_cos83;
        9'b001010100 : logcos3 = mux_in_cos84;
        9'b001010101 : logcos3 = mux_in_cos85;
        9'b001010110 : logcos3 = mux_in_cos86;
        9'b001010111 : logcos3 = mux_in_cos87;
        9'b001011000 : logcos3 = mux_in_cos88;
        9'b001011001 : logcos3 = mux_in_cos89;
        9'b001011010 : logcos3 = mux_in_cos90;
        9'b001011011 : logcos3 = mux_in_cos91;
        9'b001011100 : logcos3 = mux_in_cos92;
        9'b001011101 : logcos3 = mux_in_cos93;
        9'b001011110 : logcos3 = mux_in_cos94;
        9'b001011111 : logcos3 = mux_in_cos95;
        9'b001100000 : logcos3 = mux_in_cos96;
        9'b001100001 : logcos3 = mux_in_cos97;
        9'b001100010 : logcos3 = mux_in_cos98;
        9'b001100011 : logcos3 = mux_in_cos99;
        9'b001100100 : logcos3 = mux_in_cos100;
        9'b001100101 : logcos3 = mux_in_cos101;
        9'b001100110 : logcos3 = mux_in_cos102;
        9'b001100111 : logcos3 = mux_in_cos103;
        9'b001101000 : logcos3 = mux_in_cos104;
        9'b001101001 : logcos3 = mux_in_cos105;
        9'b001101010 : logcos3 = mux_in_cos106;
        9'b001101011 : logcos3 = mux_in_cos107;
        9'b001101100 : logcos3 = mux_in_cos108;
        9'b001101101 : logcos3 = mux_in_cos109;
        9'b001101110 : logcos3 = mux_in_cos110;
        9'b001101111 : logcos3 = mux_in_cos111;
        9'b001110000 : logcos3 = mux_in_cos112;
        9'b001110001 : logcos3 = mux_in_cos113;
        9'b001110010 : logcos3 = mux_in_cos114;
        9'b001110011 : logcos3 = mux_in_cos115;
        9'b001110100 : logcos3 = mux_in_cos116;
        9'b001110101 : logcos3 = mux_in_cos117;
        9'b001110110 : logcos3 = mux_in_cos118;
        9'b001110111 : logcos3 = mux_in_cos119;
        9'b001111000 : logcos3 = mux_in_cos120;
        9'b001111001 : logcos3 = mux_in_cos121;
        9'b001111010 : logcos3 = mux_in_cos122;
        9'b001111011 : logcos3 = mux_in_cos123;
        9'b001111100 : logcos3 = mux_in_cos124;
        9'b001111101 : logcos3 = mux_in_cos125;
        9'b001111110 : logcos3 = mux_in_cos126;
        9'b001111111 : logcos3 = mux_in_cos127;
        9'b010000000 : logcos3 = mux_in_cos128;
        9'b010000001 : logcos3 = mux_in_cos129;
        9'b010000010 : logcos3 = mux_in_cos130;
        9'b010000011 : logcos3 = mux_in_cos131;
        9'b010000100 : logcos3 = mux_in_cos132;
        9'b010000101 : logcos3 = mux_in_cos133;
        9'b010000110 : logcos3 = mux_in_cos134;
        9'b010000111 : logcos3 = mux_in_cos135;
        9'b010001000 : logcos3 = mux_in_cos136;
        9'b010001001 : logcos3 = mux_in_cos137;
        9'b010001010 : logcos3 = mux_in_cos138;
        9'b010001011 : logcos3 = mux_in_cos139;
        9'b010001100 : logcos3 = mux_in_cos140;
        9'b010001101 : logcos3 = mux_in_cos141;
        9'b010001110 : logcos3 = mux_in_cos142;
        9'b010001111 : logcos3 = mux_in_cos143;
        9'b010010000 : logcos3 = mux_in_cos144;
        9'b010010001 : logcos3 = mux_in_cos145;
        9'b010010010 : logcos3 = mux_in_cos146;
        9'b010010011 : logcos3 = mux_in_cos147;
        9'b010010100 : logcos3 = mux_in_cos148;
        9'b010010101 : logcos3 = mux_in_cos149;
        9'b010010110 : logcos3 = mux_in_cos150;
        9'b010010111 : logcos3 = mux_in_cos151;
        9'b010011000 : logcos3 = mux_in_cos152;
        9'b010011001 : logcos3 = mux_in_cos153;
        9'b010011010 : logcos3 = mux_in_cos154;
        9'b010011011 : logcos3 = mux_in_cos155;
        9'b010011100 : logcos3 = mux_in_cos156;
        9'b010011101 : logcos3 = mux_in_cos157;
        9'b010011110 : logcos3 = mux_in_cos158;
        9'b010011111 : logcos3 = mux_in_cos159;
        9'b010100000 : logcos3 = mux_in_cos160;
        9'b010100001 : logcos3 = mux_in_cos161;
        9'b010100010 : logcos3 = mux_in_cos162;
        9'b010100011 : logcos3 = mux_in_cos163;
        9'b010100100 : logcos3 = mux_in_cos164;
        9'b010100101 : logcos3 = mux_in_cos165;
        9'b010100110 : logcos3 = mux_in_cos166;
        9'b010100111 : logcos3 = mux_in_cos167;
        9'b010101000 : logcos3 = mux_in_cos168;
        9'b010101001 : logcos3 = mux_in_cos169;
        9'b010101010 : logcos3 = mux_in_cos170;
        9'b010101011 : logcos3 = mux_in_cos171;
        9'b010101100 : logcos3 = mux_in_cos172;
        9'b010101101 : logcos3 = mux_in_cos173;
        9'b010101110 : logcos3 = mux_in_cos174;
        9'b010101111 : logcos3 = mux_in_cos175;
        9'b010110000 : logcos3 = mux_in_cos176;
        9'b010110001 : logcos3 = mux_in_cos177;
        9'b010110010 : logcos3 = mux_in_cos178;
        9'b010110011 : logcos3 = mux_in_cos179;
        9'b010110100 : logcos3 = mux_in_cos180;
        9'b010110101 : logcos3 = mux_in_cos181;
        9'b010110110 : logcos3 = mux_in_cos182;
        9'b010110111 : logcos3 = mux_in_cos183;
        9'b010111000 : logcos3 = mux_in_cos184;
        9'b010111001 : logcos3 = mux_in_cos185;
        9'b010111010 : logcos3 = mux_in_cos186;
        9'b010111011 : logcos3 = mux_in_cos187;
        9'b010111100 : logcos3 = mux_in_cos188;
        9'b010111101 : logcos3 = mux_in_cos189;
        9'b010111110 : logcos3 = mux_in_cos190;
        9'b010111111 : logcos3 = mux_in_cos191;
        9'b011000000 : logcos3 = mux_in_cos192;
        9'b011000001 : logcos3 = mux_in_cos193;
        9'b011000010 : logcos3 = mux_in_cos194;
        9'b011000011 : logcos3 = mux_in_cos195;
        9'b011000100 : logcos3 = mux_in_cos196;
        9'b011000101 : logcos3 = mux_in_cos197;
        9'b011000110 : logcos3 = mux_in_cos198;
        9'b011000111 : logcos3 = mux_in_cos199;
        9'b011001000 : logcos3 = mux_in_cos200;
        9'b011001001 : logcos3 = mux_in_cos201;
        9'b011001010 : logcos3 = mux_in_cos202;
        9'b011001011 : logcos3 = mux_in_cos203;
        9'b011001100 : logcos3 = mux_in_cos204;
        9'b011001101 : logcos3 = mux_in_cos205;
        9'b011001110 : logcos3 = mux_in_cos206;
        9'b011001111 : logcos3 = mux_in_cos207;
        9'b011010000 : logcos3 = mux_in_cos208;
        9'b011010001 : logcos3 = mux_in_cos209;
        9'b011010010 : logcos3 = mux_in_cos210;
        9'b011010011 : logcos3 = mux_in_cos211;
        9'b011010100 : logcos3 = mux_in_cos212;
        9'b011010101 : logcos3 = mux_in_cos213;
        9'b011010110 : logcos3 = mux_in_cos214;
        9'b011010111 : logcos3 = mux_in_cos215;
        9'b011011000 : logcos3 = mux_in_cos216;
        9'b011011001 : logcos3 = mux_in_cos217;
        9'b011011010 : logcos3 = mux_in_cos218;
        9'b011011011 : logcos3 = mux_in_cos219;
        9'b011011100 : logcos3 = mux_in_cos220;
        9'b011011101 : logcos3 = mux_in_cos221;
        9'b011011110 : logcos3 = mux_in_cos222;
        9'b011011111 : logcos3 = mux_in_cos223;
        9'b011100000 : logcos3 = mux_in_cos224;
        9'b011100001 : logcos3 = mux_in_cos225;
        9'b011100010 : logcos3 = mux_in_cos226;
        9'b011100011 : logcos3 = mux_in_cos227;
        9'b011100100 : logcos3 = mux_in_cos228;
        9'b011100101 : logcos3 = mux_in_cos229;
        9'b011100110 : logcos3 = mux_in_cos230;
        9'b011100111 : logcos3 = mux_in_cos231;
        9'b011101000 : logcos3 = mux_in_cos232;
        9'b011101001 : logcos3 = mux_in_cos233;
        9'b011101010 : logcos3 = mux_in_cos234;
        9'b011101011 : logcos3 = mux_in_cos235;
        9'b011101100 : logcos3 = mux_in_cos236;
        9'b011101101 : logcos3 = mux_in_cos237;
        9'b011101110 : logcos3 = mux_in_cos238;
        9'b011101111 : logcos3 = mux_in_cos239;
        9'b011110000 : logcos3 = mux_in_cos240;
        9'b011110001 : logcos3 = mux_in_cos241;
        9'b011110010 : logcos3 = mux_in_cos242;
        9'b011110011 : logcos3 = mux_in_cos243;
        9'b011110100 : logcos3 = mux_in_cos244;
        9'b011110101 : logcos3 = mux_in_cos245;
        9'b011110110 : logcos3 = mux_in_cos246;
        9'b011110111 : logcos3 = mux_in_cos247;
        9'b011111000 : logcos3 = mux_in_cos248;
        9'b011111001 : logcos3 = mux_in_cos249;
        9'b011111010 : logcos3 = mux_in_cos250;
        9'b011111011 : logcos3 = mux_in_cos251;
        9'b011111100 : logcos3 = mux_in_cos252;
        9'b011111101 : logcos3 = mux_in_cos253;
        9'b011111110 : logcos3 = mux_in_cos254;
        9'b011111111 : logcos3 = mux_in_cos255;
        9'b100000000 : logcos3 = mux_in_cos256;
        default: logcos3 = 15'bx;
        endcase
    end
    
endmodule